//`include "/eda/ams/verilog/c35b3/c35_CORELIB.v"
//`include "/eda/ams/verilog/udp.v"


module Multipliers_DW_mult_tc_0 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n513, n514, n515,
         n516, n517, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1517, n1518, n1519, n1520, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562;

  ADD32 U243 ( .A(n514), .B(n515), .CI(n452), .CO(n451), .S(product[60]) );
  ADD32 U244 ( .A(n519), .B(n516), .CI(n453), .CO(n452), .S(product[59]) );
  ADD32 U245 ( .A(n523), .B(n520), .CI(n454), .CO(n453), .S(product[58]) );
  ADD32 U246 ( .A(n529), .B(n524), .CI(n455), .CO(n454), .S(product[57]) );
  ADD32 U247 ( .A(n535), .B(n530), .CI(n456), .CO(n455), .S(product[56]) );
  ADD32 U248 ( .A(n536), .B(n543), .CI(n457), .CO(n456), .S(product[55]) );
  ADD32 U249 ( .A(n544), .B(n551), .CI(n458), .CO(n457), .S(product[54]) );
  ADD32 U253 ( .A(n584), .B(n595), .CI(n462), .CO(n461), .S(product[50]) );
  ADD32 U254 ( .A(n596), .B(n609), .CI(n463), .CO(n462), .S(product[49]) );
  ADD32 U255 ( .A(n610), .B(n623), .CI(n464), .CO(n463), .S(product[48]) );
  ADD32 U256 ( .A(n624), .B(n639), .CI(n465), .CO(n464), .S(product[47]) );
  ADD32 U257 ( .A(n640), .B(n655), .CI(n466), .CO(n465), .S(product[46]) );
  ADD32 U258 ( .A(n656), .B(n673), .CI(n467), .CO(n466), .S(product[45]) );
  ADD32 U259 ( .A(n674), .B(n691), .CI(n468), .CO(n467), .S(product[44]) );
  ADD32 U263 ( .A(n754), .B(n775), .CI(n472), .CO(n471), .S(product[40]) );
  ADD32 U264 ( .A(n776), .B(n799), .CI(n473), .CO(n472), .S(product[39]) );
  ADD32 U265 ( .A(n800), .B(n823), .CI(n474), .CO(n473), .S(product[38]) );
  ADD32 U266 ( .A(n824), .B(n849), .CI(n475), .CO(n474), .S(product[37]) );
  ADD32 U267 ( .A(n850), .B(n875), .CI(n476), .CO(n475), .S(product[36]) );
  ADD32 U268 ( .A(n876), .B(n903), .CI(n477), .CO(n476), .S(product[35]) );
  ADD32 U269 ( .A(n904), .B(n931), .CI(n478), .CO(n477), .S(product[34]) );
  ADD32 U273 ( .A(n1022), .B(n1049), .CI(n482), .CO(n481), .S(product[30]) );
  ADD32 U274 ( .A(n1050), .B(n1077), .CI(n483), .CO(n482), .S(product[29]) );
  ADD32 U275 ( .A(n1078), .B(n1103), .CI(n484), .CO(n483), .S(product[28]) );
  ADD32 U276 ( .A(n1104), .B(n1129), .CI(n485), .CO(n484), .S(product[27]) );
  ADD32 U277 ( .A(n1130), .B(n1153), .CI(n486), .CO(n485), .S(product[26]) );
  ADD32 U278 ( .A(n1154), .B(n1177), .CI(n487), .CO(n486), .S(product[25]) );
  ADD32 U279 ( .A(n1178), .B(n1199), .CI(n488), .CO(n487), .S(product[24]) );
  ADD32 U283 ( .A(n1262), .B(n1279), .CI(n492), .CO(n491), .S(product[20]) );
  ADD32 U284 ( .A(n1280), .B(n1297), .CI(n493), .CO(n492), .S(product[19]) );
  ADD32 U285 ( .A(n1298), .B(n1313), .CI(n494), .CO(n493), .S(product[18]) );
  ADD32 U286 ( .A(n1314), .B(n1329), .CI(n495), .CO(n494), .S(product[17]) );
  ADD32 U287 ( .A(n1330), .B(n1343), .CI(n496), .CO(n495), .S(product[16]) );
  ADD32 U288 ( .A(n1344), .B(n1357), .CI(n497), .CO(n496), .S(product[15]) );
  ADD32 U289 ( .A(n1358), .B(n1369), .CI(n498), .CO(n497), .S(product[14]) );
  ADD32 U290 ( .A(n1370), .B(n1381), .CI(n499), .CO(n498), .S(product[13]) );
  ADD32 U291 ( .A(n1382), .B(n1391), .CI(n500), .CO(n499), .S(product[12]) );
  ADD32 U292 ( .A(n1392), .B(n1401), .CI(n501), .CO(n500), .S(product[11]) );
  ADD32 U297 ( .A(n1430), .B(n1433), .CI(n506), .CO(n505), .S(product[6]) );
  ADD32 U298 ( .A(n1434), .B(n1436), .CI(n507), .CO(n506), .S(product[5]) );
  ADD32 U299 ( .A(n1438), .B(n1439), .CI(n508), .CO(n507), .S(product[4]) );
  ADD32 U301 ( .A(n1936), .B(n1967), .CI(n510), .CO(n509), .S(product[2]) );
  ADD22 U302 ( .A(n1968), .B(n1456), .CO(n510), .S(product[1]) );
  ADD32 U304 ( .A(n1458), .B(n517), .CI(n2943), .CO(n513), .S(n514) );
  ADD32 U305 ( .A(n2942), .B(n1459), .CI(n521), .CO(n515), .S(n516) );
  ADD32 U307 ( .A(n525), .B(n2946), .CI(n522), .CO(n519), .S(n520) );
  ADD32 U308 ( .A(n1490), .B(n527), .CI(n1460), .CO(n521), .S(n522) );
  ADD32 U309 ( .A(n526), .B(n533), .CI(n531), .CO(n523), .S(n524) );
  ADD32 U316 ( .A(n1461), .B(n1491), .CI(n2945), .CO(n525), .S(n526) );
  ADD32 U318 ( .A(n532), .B(n534), .CI(n537), .CO(n529), .S(n530) );
  ADD32 U319 ( .A(n2949), .B(n1522), .CI(n539), .CO(n531), .S(n532) );
  ADD32 U320 ( .A(n1492), .B(n1462), .CI(n541), .CO(n533), .S(n534) );
  ADD32 U321 ( .A(n538), .B(n547), .CI(n545), .CO(n535), .S(n536) );
  ADD32 U322 ( .A(n549), .B(n2948), .CI(n540), .CO(n537), .S(n538) );
  ADD32 U323 ( .A(n1493), .B(n1463), .CI(n1523), .CO(n539), .S(n540) );
  ADD32 U325 ( .A(n553), .B(n548), .CI(n546), .CO(n543), .S(n544) );
  ADD32 U326 ( .A(n550), .B(n557), .CI(n555), .CO(n545), .S(n546) );
  ADD32 U327 ( .A(n1524), .B(n1494), .CI(n2952), .CO(n547), .S(n548) );
  ADD32 U328 ( .A(n1554), .B(n1464), .CI(n559), .CO(n549), .S(n550) );
  ADD32 U329 ( .A(n563), .B(n556), .CI(n554), .CO(n551), .S(n552) );
  ADD32 U330 ( .A(n558), .B(n567), .CI(n565), .CO(n553), .S(n554) );
  ADD32 U331 ( .A(n2951), .B(n1525), .CI(n569), .CO(n555), .S(n556) );
  ADD32 U332 ( .A(n1555), .B(n1495), .CI(n1465), .CO(n557), .S(n558) );
  ADD32 U334 ( .A(n573), .B(n566), .CI(n564), .CO(n561), .S(n562) );
  ADD32 U335 ( .A(n570), .B(n568), .CI(n575), .CO(n563), .S(n564) );
  ADD32 U336 ( .A(n579), .B(n2955), .CI(n577), .CO(n565), .S(n566) );
  ADD32 U337 ( .A(n1496), .B(n1556), .CI(n1586), .CO(n567), .S(n568) );
  ADD32 U338 ( .A(n581), .B(n1466), .CI(n1526), .CO(n569), .S(n570) );
  ADD32 U339 ( .A(n585), .B(n576), .CI(n574), .CO(n571), .S(n572) );
  ADD32 U340 ( .A(n589), .B(n578), .CI(n587), .CO(n573), .S(n574) );
  ADD32 U341 ( .A(n591), .B(n593), .CI(n580), .CO(n575), .S(n576) );
  ADD32 U342 ( .A(n1467), .B(n1497), .CI(n2954), .CO(n577), .S(n578) );
  ADD32 U343 ( .A(n1587), .B(n1527), .CI(n1557), .CO(n579), .S(n580) );
  ADD32 U345 ( .A(n597), .B(n588), .CI(n586), .CO(n583), .S(n584) );
  ADD32 U346 ( .A(n590), .B(n601), .CI(n599), .CO(n585), .S(n586) );
  ADD32 U347 ( .A(n592), .B(n603), .CI(n594), .CO(n587), .S(n588) );
  ADD32 U348 ( .A(n2958), .B(n1558), .CI(n605), .CO(n589), .S(n590) );
  ADD32 U349 ( .A(n1528), .B(n1588), .CI(n1618), .CO(n591), .S(n592) );
  ADD32 U350 ( .A(n607), .B(n1468), .CI(n1498), .CO(n593), .S(n594) );
  ADD32 U351 ( .A(n611), .B(n600), .CI(n598), .CO(n595), .S(n596) );
  ADD32 U352 ( .A(n602), .B(n615), .CI(n613), .CO(n597), .S(n598) );
  ADD32 U353 ( .A(n606), .B(n604), .CI(n617), .CO(n599), .S(n600) );
  ADD32 U354 ( .A(n621), .B(n2957), .CI(n619), .CO(n601), .S(n602) );
  ADD32 U355 ( .A(n1469), .B(n1559), .CI(n1499), .CO(n603), .S(n604) );
  ADD32 U356 ( .A(n1619), .B(n1529), .CI(n1589), .CO(n605), .S(n606) );
  ADD32 U358 ( .A(n625), .B(n614), .CI(n612), .CO(n609), .S(n610) );
  ADD32 U359 ( .A(n616), .B(n629), .CI(n627), .CO(n611), .S(n612) );
  ADD32 U360 ( .A(n631), .B(n622), .CI(n618), .CO(n613), .S(n614) );
  ADD32 U361 ( .A(n633), .B(n635), .CI(n620), .CO(n615), .S(n616) );
  ADD32 U362 ( .A(n1650), .B(n1500), .CI(n2961), .CO(n617), .S(n618) );
  ADD32 U363 ( .A(n1560), .B(n1620), .CI(n1590), .CO(n619), .S(n620) );
  ADD32 U364 ( .A(n637), .B(n1470), .CI(n1530), .CO(n621), .S(n622) );
  ADD32 U365 ( .A(n641), .B(n628), .CI(n626), .CO(n623), .S(n624) );
  ADD32 U366 ( .A(n630), .B(n645), .CI(n643), .CO(n625), .S(n626) );
  ADD32 U367 ( .A(n647), .B(n636), .CI(n632), .CO(n627), .S(n628) );
  ADD32 U368 ( .A(n649), .B(n651), .CI(n634), .CO(n629), .S(n630) );
  ADD32 U369 ( .A(n2960), .B(n1561), .CI(n653), .CO(n631), .S(n632) );
  ADD32 U370 ( .A(n1471), .B(n1591), .CI(n1501), .CO(n633), .S(n634) );
  ADD32 U371 ( .A(n1651), .B(n1531), .CI(n1621), .CO(n635), .S(n636) );
  ADD32 U373 ( .A(n657), .B(n644), .CI(n642), .CO(n639), .S(n640) );
  ADD32 U374 ( .A(n646), .B(n661), .CI(n659), .CO(n641), .S(n642) );
  ADD32 U375 ( .A(n663), .B(n654), .CI(n648), .CO(n643), .S(n644) );
  ADD32 U376 ( .A(n650), .B(n665), .CI(n652), .CO(n645), .S(n646) );
  ADD32 U377 ( .A(n669), .B(n2964), .CI(n667), .CO(n647), .S(n648) );
  ADD32 U378 ( .A(n1622), .B(n1562), .CI(n1652), .CO(n649), .S(n650) );
  ADD32 U379 ( .A(n1502), .B(n1592), .CI(n1532), .CO(n651), .S(n652) );
  ADD32 U380 ( .A(n1682), .B(n1472), .CI(n671), .CO(n653), .S(n654) );
  ADD32 U381 ( .A(n675), .B(n660), .CI(n658), .CO(n655), .S(n656) );
  ADD32 U382 ( .A(n662), .B(n679), .CI(n677), .CO(n657), .S(n658) );
  ADD32 U383 ( .A(n681), .B(n683), .CI(n664), .CO(n659), .S(n660) );
  ADD32 U384 ( .A(n670), .B(n668), .CI(n666), .CO(n661), .S(n662) );
  ADD32 U385 ( .A(n685), .B(n689), .CI(n687), .CO(n663), .S(n664) );
  ADD32 U386 ( .A(n1653), .B(n1683), .CI(n2963), .CO(n665), .S(n666) );
  ADD32 U387 ( .A(n1593), .B(n1533), .CI(n1623), .CO(n667), .S(n668) );
  ADD32 U388 ( .A(n1473), .B(n1563), .CI(n1503), .CO(n669), .S(n670) );
  ADD32 U390 ( .A(n693), .B(n678), .CI(n676), .CO(n673), .S(n674) );
  ADD32 U391 ( .A(n680), .B(n697), .CI(n695), .CO(n675), .S(n676) );
  ADD32 U392 ( .A(n699), .B(n684), .CI(n682), .CO(n677), .S(n678) );
  ADD32 U393 ( .A(n690), .B(n688), .CI(n701), .CO(n679), .S(n680) );
  ADD32 U394 ( .A(n703), .B(n705), .CI(n686), .CO(n681), .S(n682) );
  ADD32 U395 ( .A(n2967), .B(n1684), .CI(n707), .CO(n683), .S(n684) );
  ADD32 U396 ( .A(n1654), .B(n1564), .CI(n1594), .CO(n685), .S(n686) );
  ADD32 U397 ( .A(n1534), .B(n1624), .CI(n709), .CO(n687), .S(n688) );
  ADD32 U398 ( .A(n1714), .B(n1474), .CI(n1504), .CO(n689), .S(n690) );
  ADD32 U399 ( .A(n713), .B(n696), .CI(n694), .CO(n691), .S(n692) );
  ADD32 U400 ( .A(n698), .B(n717), .CI(n715), .CO(n693), .S(n694) );
  ADD32 U401 ( .A(n719), .B(n702), .CI(n700), .CO(n695), .S(n696) );
  ADD32 U402 ( .A(n723), .B(n708), .CI(n721), .CO(n697), .S(n698) );
  ADD32 U403 ( .A(n704), .B(n725), .CI(n706), .CO(n699), .S(n700) );
  ADD32 U404 ( .A(n729), .B(n2966), .CI(n727), .CO(n701), .S(n702) );
  ADD32 U405 ( .A(n1535), .B(n1625), .CI(n1595), .CO(n703), .S(n704) );
  ADD32 U406 ( .A(n1655), .B(n1475), .CI(n1505), .CO(n705), .S(n706) );
  ADD32 U407 ( .A(n1715), .B(n1565), .CI(n1685), .CO(n707), .S(n708) );
  ADD32 U409 ( .A(n733), .B(n716), .CI(n714), .CO(n711), .S(n712) );
  ADD32 U410 ( .A(n718), .B(n737), .CI(n735), .CO(n713), .S(n714) );
  ADD32 U411 ( .A(n722), .B(n739), .CI(n720), .CO(n715), .S(n716) );
  ADD32 U412 ( .A(n741), .B(n743), .CI(n724), .CO(n717), .S(n718) );
  ADD32 U413 ( .A(n730), .B(n726), .CI(n728), .CO(n719), .S(n720) );
  ADD32 U414 ( .A(n745), .B(n749), .CI(n747), .CO(n721), .S(n722) );
  ADD32 U415 ( .A(n1686), .B(n1716), .CI(n2970), .CO(n723), .S(n724) );
  ADD32 U416 ( .A(n1656), .B(n1536), .CI(n1596), .CO(n725), .S(n726) );
  ADD32 U417 ( .A(n751), .B(n1626), .CI(n1566), .CO(n727), .S(n728) );
  ADD32 U418 ( .A(n1746), .B(n1476), .CI(n1506), .CO(n729), .S(n730) );
  ADD32 U419 ( .A(n755), .B(n736), .CI(n734), .CO(n731), .S(n732) );
  ADD32 U420 ( .A(n738), .B(n759), .CI(n757), .CO(n733), .S(n734) );
  ADD32 U421 ( .A(n742), .B(n761), .CI(n740), .CO(n735), .S(n736) );
  ADD32 U422 ( .A(n744), .B(n765), .CI(n763), .CO(n737), .S(n738) );
  ADD32 U423 ( .A(n750), .B(n746), .CI(n748), .CO(n739), .S(n740) );
  ADD32 U424 ( .A(n767), .B(n771), .CI(n769), .CO(n741), .S(n742) );
  ADD32 U425 ( .A(n2969), .B(n1657), .CI(n773), .CO(n743), .S(n744) );
  ADD32 U426 ( .A(n1537), .B(n1687), .CI(n1627), .CO(n745), .S(n746) );
  ADD32 U427 ( .A(n1507), .B(n1567), .CI(n1717), .CO(n747), .S(n748) );
  ADD32 U428 ( .A(n1477), .B(n1597), .CI(n1747), .CO(n749), .S(n750) );
  ADD32 U430 ( .A(n777), .B(n758), .CI(n756), .CO(n753), .S(n754) );
  ADD32 U431 ( .A(n760), .B(n781), .CI(n779), .CO(n755), .S(n756) );
  ADD32 U432 ( .A(n783), .B(n764), .CI(n762), .CO(n757), .S(n758) );
  ADD32 U433 ( .A(n766), .B(n787), .CI(n785), .CO(n759), .S(n760) );
  ADD32 U434 ( .A(n774), .B(n770), .CI(n772), .CO(n761), .S(n762) );
  ADD32 U435 ( .A(n789), .B(n791), .CI(n768), .CO(n763), .S(n764) );
  ADD32 U436 ( .A(n795), .B(n2973), .CI(n793), .CO(n765), .S(n766) );
  ADD32 U437 ( .A(n1628), .B(n1778), .CI(n1748), .CO(n767), .S(n768) );
  ADD32 U438 ( .A(n1598), .B(n1658), .CI(n1718), .CO(n769), .S(n770) );
  ADD32 U439 ( .A(n1568), .B(n1688), .CI(n1508), .CO(n771), .S(n772) );
  ADD32 U440 ( .A(n797), .B(n1478), .CI(n1538), .CO(n773), .S(n774) );
  ADD32 U441 ( .A(n801), .B(n780), .CI(n778), .CO(n775), .S(n776) );
  ADD32 U442 ( .A(n782), .B(n805), .CI(n803), .CO(n777), .S(n778) );
  ADD32 U443 ( .A(n807), .B(n786), .CI(n784), .CO(n779), .S(n780) );
  ADD32 U444 ( .A(n809), .B(n811), .CI(n788), .CO(n781), .S(n782) );
  ADD32 U445 ( .A(n790), .B(n796), .CI(n813), .CO(n783), .S(n784) );
  ADD32 U446 ( .A(n792), .B(n819), .CI(n794), .CO(n785), .S(n786) );
  ADD32 U447 ( .A(n815), .B(n821), .CI(n817), .CO(n787), .S(n788) );
  ADD32 U448 ( .A(n1599), .B(n1689), .CI(n2972), .CO(n789), .S(n790) );
  ADD32 U449 ( .A(n1539), .B(n1719), .CI(n1569), .CO(n791), .S(n792) );
  ADD32 U450 ( .A(n1779), .B(n1659), .CI(n1749), .CO(n793), .S(n794) );
  ADD32 U451 ( .A(n1479), .B(n1629), .CI(n1509), .CO(n795), .S(n796) );
  ADD32 U453 ( .A(n825), .B(n804), .CI(n802), .CO(n799), .S(n800) );
  ADD32 U454 ( .A(n806), .B(n829), .CI(n827), .CO(n801), .S(n802) );
  ADD32 U455 ( .A(n831), .B(n810), .CI(n808), .CO(n803), .S(n804) );
  ADD32 U456 ( .A(n833), .B(n835), .CI(n812), .CO(n805), .S(n806) );
  ADD32 U457 ( .A(n837), .B(n818), .CI(n814), .CO(n807), .S(n808) );
  ADD32 U458 ( .A(n822), .B(n816), .CI(n820), .CO(n809), .S(n810) );
  ADD32 U459 ( .A(n841), .B(n839), .CI(n843), .CO(n811), .S(n812) );
  ADD32 U460 ( .A(n2976), .B(n1780), .CI(n845), .CO(n813), .S(n814) );
  ADD32 U461 ( .A(n1510), .B(n1750), .CI(n1720), .CO(n815), .S(n816) );
  ADD32 U462 ( .A(n1600), .B(n1690), .CI(n1630), .CO(n817), .S(n818) );
  ADD32 U463 ( .A(n1540), .B(n1660), .CI(n1570), .CO(n819), .S(n820) );
  ADD32 U464 ( .A(n1810), .B(n1480), .CI(n847), .CO(n821), .S(n822) );
  ADD32 U465 ( .A(n851), .B(n828), .CI(n826), .CO(n823), .S(n824) );
  ADD32 U466 ( .A(n830), .B(n855), .CI(n853), .CO(n825), .S(n826) );
  ADD32 U467 ( .A(n857), .B(n834), .CI(n832), .CO(n827), .S(n828) );
  ADD32 U468 ( .A(n836), .B(n861), .CI(n859), .CO(n829), .S(n830) );
  ADD32 U469 ( .A(n863), .B(n865), .CI(n838), .CO(n831), .S(n832) );
  ADD32 U470 ( .A(n846), .B(n842), .CI(n844), .CO(n833), .S(n834) );
  ADD32 U471 ( .A(n867), .B(n869), .CI(n840), .CO(n835), .S(n836) );
  ADD32 U472 ( .A(n873), .B(n2975), .CI(n871), .CO(n837), .S(n838) );
  ADD32 U473 ( .A(n1661), .B(n1721), .CI(n1691), .CO(n839), .S(n840) );
  ADD32 U474 ( .A(n1541), .B(n1751), .CI(n1601), .CO(n841), .S(n842) );
  ADD32 U475 ( .A(n1481), .B(n1571), .CI(n1511), .CO(n843), .S(n844) );
  ADD32 U476 ( .A(n1811), .B(n1631), .CI(n1781), .CO(n845), .S(n846) );
  ADD32 U478 ( .A(n877), .B(n854), .CI(n852), .CO(n849), .S(n850) );
  ADD32 U479 ( .A(n856), .B(n881), .CI(n879), .CO(n851), .S(n852) );
  ADD32 U480 ( .A(n883), .B(n860), .CI(n858), .CO(n853), .S(n854) );
  ADD32 U481 ( .A(n885), .B(n864), .CI(n862), .CO(n855), .S(n856) );
  ADD32 U482 ( .A(n866), .B(n889), .CI(n887), .CO(n857), .S(n858) );
  ADD32 U483 ( .A(n874), .B(n872), .CI(n891), .CO(n859), .S(n860) );
  ADD32 U484 ( .A(n868), .B(n897), .CI(n870), .CO(n861), .S(n862) );
  ADD32 U485 ( .A(n899), .B(n895), .CI(n893), .CO(n863), .S(n864) );
  ADD32 U486 ( .A(n1782), .B(n1812), .CI(n2979), .CO(n865), .S(n866) );
  ADD32 U487 ( .A(n1752), .B(n1632), .CI(n1662), .CO(n867), .S(n868) );
  ADD32 U488 ( .A(n901), .B(n1722), .CI(n1602), .CO(n869), .S(n870) );
  ADD32 U489 ( .A(n1542), .B(n1692), .CI(n1572), .CO(n871), .S(n872) );
  ADD32 U490 ( .A(n1842), .B(n1482), .CI(n1512), .CO(n873), .S(n874) );
  ADD32 U491 ( .A(n905), .B(n880), .CI(n878), .CO(n875), .S(n876) );
  ADD32 U492 ( .A(n882), .B(n909), .CI(n907), .CO(n877), .S(n878) );
  ADD32 U493 ( .A(n911), .B(n886), .CI(n884), .CO(n879), .S(n880) );
  ADD32 U494 ( .A(n913), .B(n890), .CI(n888), .CO(n881), .S(n882) );
  ADD32 U495 ( .A(n892), .B(n917), .CI(n915), .CO(n883), .S(n884) );
  ADD32 U496 ( .A(n900), .B(n898), .CI(n919), .CO(n885), .S(n886) );
  ADD32 U497 ( .A(n894), .B(n925), .CI(n896), .CO(n887), .S(n888) );
  ADD32 U498 ( .A(n927), .B(n923), .CI(n921), .CO(n889), .S(n890) );
  ADD32 U499 ( .A(n2978), .B(n1783), .CI(n929), .CO(n891), .S(n892) );
  ADD32 U500 ( .A(n1723), .B(n1813), .CI(n1753), .CO(n893), .S(n894) );
  ADD32 U501 ( .A(n1603), .B(n1573), .CI(n1693), .CO(n895), .S(n896) );
  ADD32 U502 ( .A(n1513), .B(n1633), .CI(n1543), .CO(n897), .S(n898) );
  ADD32 U503 ( .A(n1483), .B(n1663), .CI(n1843), .CO(n899), .S(n900) );
  ADD32 U505 ( .A(n933), .B(n908), .CI(n906), .CO(n903), .S(n904) );
  ADD32 U506 ( .A(n910), .B(n937), .CI(n935), .CO(n905), .S(n906) );
  ADD32 U507 ( .A(n939), .B(n914), .CI(n912), .CO(n907), .S(n908) );
  ADD32 U508 ( .A(n941), .B(n918), .CI(n916), .CO(n909), .S(n910) );
  ADD32 U509 ( .A(n920), .B(n945), .CI(n943), .CO(n911), .S(n912) );
  ADD32 U510 ( .A(n926), .B(n924), .CI(n947), .CO(n913), .S(n914) );
  ADD32 U511 ( .A(n930), .B(n922), .CI(n928), .CO(n915), .S(n916) );
  ADD32 U512 ( .A(n951), .B(n953), .CI(n949), .CO(n917), .S(n918) );
  ADD32 U513 ( .A(n957), .B(n2982), .CI(n955), .CO(n919), .S(n920) );
  ADD32 U514 ( .A(n1874), .B(n1844), .CI(n1694), .CO(n921), .S(n922) );
  ADD32 U515 ( .A(n1784), .B(n1574), .CI(n1814), .CO(n923), .S(n924) );
  ADD32 U516 ( .A(n1634), .B(n1754), .CI(n1664), .CO(n925), .S(n926) );
  ADD32 U517 ( .A(n1544), .B(n1724), .CI(n1604), .CO(n927), .S(n928) );
  ADD32 U518 ( .A(n959), .B(n1484), .CI(n1514), .CO(n929), .S(n930) );
  ADD32 U519 ( .A(n963), .B(n936), .CI(n934), .CO(n931), .S(n932) );
  ADD32 U520 ( .A(n938), .B(n940), .CI(n965), .CO(n933), .S(n934) );
  ADD32 U521 ( .A(n969), .B(n942), .CI(n967), .CO(n935), .S(n936) );
  ADD32 U522 ( .A(n944), .B(n946), .CI(n971), .CO(n937), .S(n938) );
  ADD32 U523 ( .A(n948), .B(n975), .CI(n973), .CO(n939), .S(n940) );
  ADD32 U524 ( .A(n950), .B(n979), .CI(n977), .CO(n941), .S(n942) );
  ADD32 U525 ( .A(n958), .B(n956), .CI(n954), .CO(n943), .S(n944) );
  ADD32 U526 ( .A(n981), .B(n985), .CI(n952), .CO(n945), .S(n946) );
  ADD32 U527 ( .A(n983), .B(n2941), .CI(n987), .CO(n947), .S(n948) );
  ADD32 U528 ( .A(n1785), .B(n1755), .CI(n2981), .CO(n949), .S(n950) );
  ADD32 U529 ( .A(n1635), .B(n1815), .CI(n1725), .CO(n951), .S(n952) );
  ADD32 U530 ( .A(n1845), .B(n1575), .CI(n1605), .CO(n953), .S(n954) );
  ADD32 U531 ( .A(n1875), .B(n1695), .CI(n1545), .CO(n955), .S(n956) );
  ADD32 U532 ( .A(n1485), .B(n1665), .CI(n1515), .CO(n957), .S(n958) );
  ADD32 U534 ( .A(n993), .B(n966), .CI(n964), .CO(n961), .S(n962) );
  ADD32 U535 ( .A(n968), .B(n970), .CI(n995), .CO(n963), .S(n964) );
  ADD32 U536 ( .A(n999), .B(n972), .CI(n997), .CO(n965), .S(n966) );
  ADD32 U537 ( .A(n1001), .B(n976), .CI(n974), .CO(n967), .S(n968) );
  ADD32 U538 ( .A(n1003), .B(n980), .CI(n978), .CO(n969), .S(n970) );
  ADD32 U539 ( .A(n1007), .B(n990), .CI(n1005), .CO(n971), .S(n972) );
  ADD32 U540 ( .A(n988), .B(n984), .CI(n986), .CO(n973), .S(n974) );
  ADD32 U541 ( .A(n1013), .B(n1009), .CI(n982), .CO(n975), .S(n976) );
  ADD32 U542 ( .A(n1017), .B(n1011), .CI(n1015), .CO(n977), .S(n978) );
  ADD32 U543 ( .A(n2984), .B(n1846), .CI(n1019), .CO(n979), .S(n980) );
  ADD32 U544 ( .A(n1816), .B(n1876), .CI(n1906), .CO(n981), .S(n982) );
  ADD32 U545 ( .A(n1636), .B(n1726), .CI(n1666), .CO(n983), .S(n984) );
  ADD32 U546 ( .A(n1606), .B(n1786), .CI(n1576), .CO(n985), .S(n986) );
  ADD32 U547 ( .A(n1546), .B(n1696), .CI(n1486), .CO(n987), .S(n988) );
  ADD32 U549 ( .A(n1023), .B(n996), .CI(n994), .CO(n991), .S(n992) );
  ADD32 U550 ( .A(n998), .B(n1000), .CI(n1025), .CO(n993), .S(n994) );
  ADD32 U551 ( .A(n1029), .B(n1002), .CI(n1027), .CO(n995), .S(n996) );
  ADD32 U552 ( .A(n1031), .B(n1006), .CI(n1004), .CO(n997), .S(n998) );
  ADD32 U553 ( .A(n1033), .B(n1035), .CI(n1008), .CO(n999), .S(n1000) );
  ADD32 U554 ( .A(n1014), .B(n1012), .CI(n1037), .CO(n1001), .S(n1002) );
  ADD32 U555 ( .A(n1018), .B(n1010), .CI(n1016), .CO(n1003), .S(n1004) );
  ADD32 U556 ( .A(n1043), .B(n1020), .CI(n1039), .CO(n1005), .S(n1006) );
  ADD32 U557 ( .A(n1045), .B(n1047), .CI(n1041), .CO(n1007), .S(n1008) );
  ADD32 U558 ( .A(n1727), .B(n1607), .CI(n1667), .CO(n1009), .S(n1010) );
  ADD32 U559 ( .A(n1547), .B(n1757), .CI(n1577), .CO(n1011), .S(n1012) );
  ADD32 U560 ( .A(n1817), .B(n1637), .CI(n1787), .CO(n1013), .S(n1014) );
  ADD32 U561 ( .A(n1877), .B(n1697), .CI(n1847), .CO(n1015), .S(n1016) );
  ADD32 U562 ( .A(n1487), .B(n1907), .CI(n1517), .CO(n1017), .S(n1018) );
  ADD22 U563 ( .A(n1441), .B(n1938), .CO(n1019), .S(n1020) );
  ADD32 U564 ( .A(n1051), .B(n1026), .CI(n1024), .CO(n1021), .S(n1022) );
  ADD32 U565 ( .A(n1028), .B(n1030), .CI(n1053), .CO(n1023), .S(n1024) );
  ADD32 U566 ( .A(n1057), .B(n1032), .CI(n1055), .CO(n1025), .S(n1026) );
  ADD32 U567 ( .A(n1036), .B(n1059), .CI(n1034), .CO(n1027), .S(n1028) );
  ADD32 U568 ( .A(n1038), .B(n1063), .CI(n1061), .CO(n1029), .S(n1030) );
  ADD32 U569 ( .A(n1040), .B(n1042), .CI(n1065), .CO(n1031), .S(n1032) );
  ADD32 U570 ( .A(n1046), .B(n1048), .CI(n1044), .CO(n1033), .S(n1034) );
  ADD32 U571 ( .A(n1073), .B(n1069), .CI(n1071), .CO(n1035), .S(n1036) );
  ADD32 U572 ( .A(n1075), .B(n1788), .CI(n1067), .CO(n1037), .S(n1038) );
  ADD32 U573 ( .A(n1728), .B(n1818), .CI(n1758), .CO(n1039), .S(n1040) );
  ADD32 U574 ( .A(n1668), .B(n1638), .CI(n1698), .CO(n1041), .S(n1042) );
  ADD32 U575 ( .A(n1578), .B(n1848), .CI(n1608), .CO(n1043), .S(n1044) );
  ADD32 U576 ( .A(n1548), .B(n1878), .CI(n1488), .CO(n1045), .S(n1046) );
  ADD32 U577 ( .A(n1908), .B(n1939), .CI(n1518), .CO(n1047), .S(n1048) );
  ADD32 U578 ( .A(n1079), .B(n1054), .CI(n1052), .CO(n1049), .S(n1050) );
  ADD32 U579 ( .A(n1056), .B(n1058), .CI(n1081), .CO(n1051), .S(n1052) );
  ADD32 U580 ( .A(n1085), .B(n1060), .CI(n1083), .CO(n1053), .S(n1054) );
  ADD32 U581 ( .A(n1087), .B(n1064), .CI(n1062), .CO(n1055), .S(n1056) );
  ADD32 U582 ( .A(n1066), .B(n1091), .CI(n1089), .CO(n1057), .S(n1058) );
  ADD32 U583 ( .A(n1070), .B(n1072), .CI(n1074), .CO(n1059), .S(n1060) );
  ADD32 U584 ( .A(n1093), .B(n1095), .CI(n1068), .CO(n1061), .S(n1062) );
  ADD32 U585 ( .A(n1099), .B(n1076), .CI(n1097), .CO(n1063), .S(n1064) );
  ADD32 U586 ( .A(n1759), .B(n1729), .CI(n1101), .CO(n1065), .S(n1066) );
  ADD32 U587 ( .A(n1639), .B(n1789), .CI(n1699), .CO(n1067), .S(n1068) );
  ADD32 U588 ( .A(n1549), .B(n1609), .CI(n1579), .CO(n1069), .S(n1070) );
  ADD32 U589 ( .A(n1849), .B(n1669), .CI(n1819), .CO(n1071), .S(n1072) );
  ADD32 U590 ( .A(n1519), .B(n1909), .CI(n1879), .CO(n1073), .S(n1074) );
  ADD22 U591 ( .A(n1442), .B(n1940), .CO(n1075), .S(n1076) );
  ADD32 U592 ( .A(n1105), .B(n1082), .CI(n1080), .CO(n1077), .S(n1078) );
  ADD32 U593 ( .A(n1084), .B(n1109), .CI(n1107), .CO(n1079), .S(n1080) );
  ADD32 U594 ( .A(n1088), .B(n1111), .CI(n1086), .CO(n1081), .S(n1082) );
  ADD32 U595 ( .A(n1113), .B(n1092), .CI(n1090), .CO(n1083), .S(n1084) );
  ADD32 U596 ( .A(n1117), .B(n1096), .CI(n1115), .CO(n1085), .S(n1086) );
  ADD32 U597 ( .A(n1100), .B(n1094), .CI(n1098), .CO(n1087), .S(n1088) );
  ADD32 U598 ( .A(n1125), .B(n1123), .CI(n1102), .CO(n1089), .S(n1090) );
  ADD32 U599 ( .A(n1119), .B(n1127), .CI(n1121), .CO(n1091), .S(n1092) );
  ADD32 U600 ( .A(n1730), .B(n1790), .CI(n1760), .CO(n1093), .S(n1094) );
  ADD32 U601 ( .A(n1670), .B(n1820), .CI(n1700), .CO(n1095), .S(n1096) );
  ADD32 U602 ( .A(n1610), .B(n1850), .CI(n1640), .CO(n1097), .S(n1098) );
  ADD32 U603 ( .A(n1580), .B(n1880), .CI(n1520), .CO(n1099), .S(n1100) );
  ADD32 U604 ( .A(n1910), .B(n1941), .CI(n1550), .CO(n1101), .S(n1102) );
  ADD32 U605 ( .A(n1131), .B(n1108), .CI(n1106), .CO(n1103), .S(n1104) );
  ADD32 U606 ( .A(n1110), .B(n1135), .CI(n1133), .CO(n1105), .S(n1106) );
  ADD32 U607 ( .A(n1114), .B(n1137), .CI(n1112), .CO(n1107), .S(n1108) );
  ADD32 U608 ( .A(n1139), .B(n1118), .CI(n1116), .CO(n1109), .S(n1110) );
  ADD32 U609 ( .A(n1122), .B(n1124), .CI(n1141), .CO(n1111), .S(n1112) );
  ADD32 U610 ( .A(n1126), .B(n1120), .CI(n1143), .CO(n1113), .S(n1114) );
  ADD32 U611 ( .A(n1147), .B(n1145), .CI(n1149), .CO(n1115), .S(n1116) );
  ADD32 U612 ( .A(n1151), .B(n1791), .CI(n1128), .CO(n1117), .S(n1118) );
  ADD32 U613 ( .A(n1701), .B(n1821), .CI(n1761), .CO(n1119), .S(n1120) );
  ADD32 U614 ( .A(n1641), .B(n1851), .CI(n1671), .CO(n1121), .S(n1122) );
  ADD32 U615 ( .A(n1611), .B(n1731), .CI(n1881), .CO(n1123), .S(n1124) );
  ADD32 U616 ( .A(n1551), .B(n1911), .CI(n1581), .CO(n1125), .S(n1126) );
  ADD22 U617 ( .A(n1443), .B(n1942), .CO(n1127), .S(n1128) );
  ADD32 U618 ( .A(n1155), .B(n1134), .CI(n1132), .CO(n1129), .S(n1130) );
  ADD32 U619 ( .A(n1136), .B(n1159), .CI(n1157), .CO(n1131), .S(n1132) );
  ADD32 U620 ( .A(n1140), .B(n1142), .CI(n1138), .CO(n1133), .S(n1134) );
  ADD32 U621 ( .A(n1163), .B(n1144), .CI(n1161), .CO(n1135), .S(n1136) );
  ADD32 U622 ( .A(n1150), .B(n1148), .CI(n1165), .CO(n1137), .S(n1138) );
  ADD32 U623 ( .A(n1152), .B(n1171), .CI(n1146), .CO(n1139), .S(n1140) );
  ADD32 U624 ( .A(n1167), .B(n1173), .CI(n1169), .CO(n1141), .S(n1142) );
  ADD32 U625 ( .A(n1762), .B(n1792), .CI(n1175), .CO(n1143), .S(n1144) );
  ADD32 U626 ( .A(n1702), .B(n1822), .CI(n1732), .CO(n1145), .S(n1146) );
  ADD32 U627 ( .A(n1642), .B(n1852), .CI(n1672), .CO(n1147), .S(n1148) );
  ADD32 U628 ( .A(n1612), .B(n1882), .CI(n1552), .CO(n1149), .S(n1150) );
  ADD32 U629 ( .A(n1912), .B(n1943), .CI(n1582), .CO(n1151), .S(n1152) );
  ADD32 U630 ( .A(n1179), .B(n1158), .CI(n1156), .CO(n1153), .S(n1154) );
  ADD32 U631 ( .A(n1160), .B(n1183), .CI(n1181), .CO(n1155), .S(n1156) );
  ADD32 U632 ( .A(n1164), .B(n1185), .CI(n1162), .CO(n1157), .S(n1158) );
  ADD32 U633 ( .A(n1187), .B(n1189), .CI(n1166), .CO(n1159), .S(n1160) );
  ADD32 U634 ( .A(n1174), .B(n1170), .CI(n1172), .CO(n1161), .S(n1162) );
  ADD32 U635 ( .A(n1193), .B(n1176), .CI(n1168), .CO(n1163), .S(n1164) );
  ADD32 U636 ( .A(n1195), .B(n1197), .CI(n1191), .CO(n1165), .S(n1166) );
  ADD32 U637 ( .A(n1763), .B(n1823), .CI(n1793), .CO(n1167), .S(n1168) );
  ADD32 U638 ( .A(n1673), .B(n1853), .CI(n1733), .CO(n1169), .S(n1170) );
  ADD32 U639 ( .A(n1613), .B(n1703), .CI(n1643), .CO(n1171), .S(n1172) );
  ADD32 U640 ( .A(n1583), .B(n1913), .CI(n1883), .CO(n1173), .S(n1174) );
  ADD22 U641 ( .A(n1444), .B(n1944), .CO(n1175), .S(n1176) );
  ADD32 U642 ( .A(n1201), .B(n1182), .CI(n1180), .CO(n1177), .S(n1178) );
  ADD32 U643 ( .A(n1184), .B(n1205), .CI(n1203), .CO(n1179), .S(n1180) );
  ADD32 U644 ( .A(n1188), .B(n1207), .CI(n1186), .CO(n1181), .S(n1182) );
  ADD32 U645 ( .A(n1209), .B(n1211), .CI(n1190), .CO(n1183), .S(n1184) );
  ADD32 U646 ( .A(n1196), .B(n1192), .CI(n1194), .CO(n1185), .S(n1186) );
  ADD32 U647 ( .A(n1213), .B(n1215), .CI(n1198), .CO(n1187), .S(n1188) );
  ADD32 U648 ( .A(n1219), .B(n1764), .CI(n1217), .CO(n1189), .S(n1190) );
  ADD32 U649 ( .A(n1704), .B(n1794), .CI(n1734), .CO(n1191), .S(n1192) );
  ADD32 U650 ( .A(n1674), .B(n1854), .CI(n1824), .CO(n1193), .S(n1194) );
  ADD32 U651 ( .A(n1644), .B(n1884), .CI(n1584), .CO(n1195), .S(n1196) );
  ADD32 U652 ( .A(n1914), .B(n1945), .CI(n1614), .CO(n1197), .S(n1198) );
  ADD32 U653 ( .A(n1223), .B(n1204), .CI(n1202), .CO(n1199), .S(n1200) );
  ADD32 U654 ( .A(n1225), .B(n1208), .CI(n1206), .CO(n1201), .S(n1202) );
  ADD32 U655 ( .A(n1210), .B(n1229), .CI(n1227), .CO(n1203), .S(n1204) );
  ADD32 U656 ( .A(n1231), .B(n1218), .CI(n1212), .CO(n1205), .S(n1206) );
  ADD32 U657 ( .A(n1214), .B(n1237), .CI(n1216), .CO(n1207), .S(n1208) );
  ADD32 U658 ( .A(n1233), .B(n1220), .CI(n1235), .CO(n1209), .S(n1210) );
  ADD32 U659 ( .A(n1765), .B(n1795), .CI(n1239), .CO(n1211), .S(n1212) );
  ADD32 U660 ( .A(n1675), .B(n1825), .CI(n1705), .CO(n1213), .S(n1214) );
  ADD32 U661 ( .A(n1885), .B(n1735), .CI(n1855), .CO(n1215), .S(n1216) );
  ADD32 U662 ( .A(n1615), .B(n1915), .CI(n1645), .CO(n1217), .S(n1218) );
  ADD22 U663 ( .A(n1445), .B(n1946), .CO(n1219), .S(n1220) );
  ADD32 U664 ( .A(n1243), .B(n1226), .CI(n1224), .CO(n1221), .S(n1222) );
  ADD32 U665 ( .A(n1228), .B(n1230), .CI(n1245), .CO(n1223), .S(n1224) );
  ADD32 U666 ( .A(n1232), .B(n1249), .CI(n1247), .CO(n1225), .S(n1226) );
  ADD32 U667 ( .A(n1238), .B(n1236), .CI(n1251), .CO(n1227), .S(n1228) );
  ADD32 U668 ( .A(n1240), .B(n1253), .CI(n1234), .CO(n1229), .S(n1230) );
  ADD32 U669 ( .A(n1257), .B(n1259), .CI(n1255), .CO(n1231), .S(n1232) );
  ADD32 U670 ( .A(n1766), .B(n1826), .CI(n1796), .CO(n1233), .S(n1234) );
  ADD32 U671 ( .A(n1706), .B(n1856), .CI(n1736), .CO(n1235), .S(n1236) );
  ADD32 U672 ( .A(n1676), .B(n1886), .CI(n1616), .CO(n1237), .S(n1238) );
  ADD32 U673 ( .A(n1916), .B(n1947), .CI(n1646), .CO(n1239), .S(n1240) );
  ADD32 U674 ( .A(n1263), .B(n1246), .CI(n1244), .CO(n1241), .S(n1242) );
  ADD32 U675 ( .A(n1248), .B(n1250), .CI(n1265), .CO(n1243), .S(n1244) );
  ADD32 U676 ( .A(n1252), .B(n1269), .CI(n1267), .CO(n1245), .S(n1246) );
  ADD32 U677 ( .A(n1258), .B(n1256), .CI(n1271), .CO(n1247), .S(n1248) );
  ADD32 U678 ( .A(n1273), .B(n1275), .CI(n1254), .CO(n1249), .S(n1250) );
  ADD32 U679 ( .A(n1277), .B(n1767), .CI(n1260), .CO(n1251), .S(n1252) );
  ADD32 U680 ( .A(n1677), .B(n1797), .CI(n1707), .CO(n1253), .S(n1254) );
  ADD32 U681 ( .A(n1857), .B(n1737), .CI(n1827), .CO(n1255), .S(n1256) );
  ADD32 U682 ( .A(n1647), .B(n1917), .CI(n1887), .CO(n1257), .S(n1258) );
  ADD22 U683 ( .A(n1446), .B(n1948), .CO(n1259), .S(n1260) );
  ADD32 U684 ( .A(n1281), .B(n1266), .CI(n1264), .CO(n1261), .S(n1262) );
  ADD32 U685 ( .A(n1268), .B(n1270), .CI(n1283), .CO(n1263), .S(n1264) );
  ADD32 U686 ( .A(n1272), .B(n1287), .CI(n1285), .CO(n1265), .S(n1266) );
  ADD32 U687 ( .A(n1276), .B(n1278), .CI(n1274), .CO(n1267), .S(n1268) );
  ADD32 U688 ( .A(n1289), .B(n1293), .CI(n1291), .CO(n1269), .S(n1270) );
  ADD32 U689 ( .A(n1798), .B(n1828), .CI(n1295), .CO(n1271), .S(n1272) );
  ADD32 U690 ( .A(n1738), .B(n1858), .CI(n1768), .CO(n1273), .S(n1274) );
  ADD32 U691 ( .A(n1708), .B(n1888), .CI(n1648), .CO(n1275), .S(n1276) );
  ADD32 U692 ( .A(n1918), .B(n1949), .CI(n1678), .CO(n1277), .S(n1278) );
  ADD32 U693 ( .A(n1299), .B(n1284), .CI(n1282), .CO(n1279), .S(n1280) );
  ADD32 U694 ( .A(n1286), .B(n1288), .CI(n1301), .CO(n1281), .S(n1282) );
  ADD32 U695 ( .A(n1305), .B(n1294), .CI(n1303), .CO(n1283), .S(n1284) );
  ADD32 U696 ( .A(n1290), .B(n1296), .CI(n1292), .CO(n1285), .S(n1286) );
  ADD32 U697 ( .A(n1309), .B(n1311), .CI(n1307), .CO(n1287), .S(n1288) );
  ADD32 U698 ( .A(n1769), .B(n1859), .CI(n1829), .CO(n1289), .S(n1290) );
  ADD32 U699 ( .A(n1889), .B(n1799), .CI(n1739), .CO(n1291), .S(n1292) );
  ADD32 U700 ( .A(n1679), .B(n1919), .CI(n1709), .CO(n1293), .S(n1294) );
  ADD22 U701 ( .A(n1447), .B(n1950), .CO(n1295), .S(n1296) );
  ADD32 U702 ( .A(n1315), .B(n1302), .CI(n1300), .CO(n1297), .S(n1298) );
  ADD32 U703 ( .A(n1304), .B(n1306), .CI(n1317), .CO(n1299), .S(n1300) );
  ADD32 U704 ( .A(n1321), .B(n1310), .CI(n1319), .CO(n1301), .S(n1302) );
  ADD32 U705 ( .A(n1312), .B(n1323), .CI(n1308), .CO(n1303), .S(n1304) );
  ADD32 U706 ( .A(n1327), .B(n1830), .CI(n1325), .CO(n1305), .S(n1306) );
  ADD32 U707 ( .A(n1770), .B(n1860), .CI(n1800), .CO(n1307), .S(n1308) );
  ADD32 U708 ( .A(n1740), .B(n1890), .CI(n1680), .CO(n1309), .S(n1310) );
  ADD32 U709 ( .A(n1920), .B(n1951), .CI(n1710), .CO(n1311), .S(n1312) );
  ADD32 U710 ( .A(n1331), .B(n1318), .CI(n1316), .CO(n1313), .S(n1314) );
  ADD32 U711 ( .A(n1333), .B(n1322), .CI(n1320), .CO(n1315), .S(n1316) );
  ADD32 U712 ( .A(n1326), .B(n1324), .CI(n1335), .CO(n1317), .S(n1318) );
  ADD32 U713 ( .A(n1337), .B(n1328), .CI(n1339), .CO(n1319), .S(n1320) );
  ADD32 U714 ( .A(n1831), .B(n1861), .CI(n1341), .CO(n1321), .S(n1322) );
  ADD32 U715 ( .A(n1741), .B(n1771), .CI(n1801), .CO(n1323), .S(n1324) );
  ADD32 U716 ( .A(n1711), .B(n1921), .CI(n1891), .CO(n1325), .S(n1326) );
  ADD22 U717 ( .A(n1448), .B(n1952), .CO(n1327), .S(n1328) );
  ADD32 U718 ( .A(n1345), .B(n1334), .CI(n1332), .CO(n1329), .S(n1330) );
  ADD32 U719 ( .A(n1336), .B(n1349), .CI(n1347), .CO(n1331), .S(n1332) );
  ADD32 U720 ( .A(n1340), .B(n1342), .CI(n1338), .CO(n1333), .S(n1334) );
  ADD32 U721 ( .A(n1353), .B(n1355), .CI(n1351), .CO(n1335), .S(n1336) );
  ADD32 U722 ( .A(n1802), .B(n1862), .CI(n1832), .CO(n1337), .S(n1338) );
  ADD32 U723 ( .A(n1772), .B(n1892), .CI(n1712), .CO(n1339), .S(n1340) );
  ADD32 U724 ( .A(n1922), .B(n1953), .CI(n1742), .CO(n1341), .S(n1342) );
  ADD32 U725 ( .A(n1359), .B(n1348), .CI(n1346), .CO(n1343), .S(n1344) );
  ADD32 U726 ( .A(n1361), .B(n1363), .CI(n1350), .CO(n1345), .S(n1346) );
  ADD32 U727 ( .A(n1352), .B(n1365), .CI(n1354), .CO(n1347), .S(n1348) );
  ADD32 U728 ( .A(n1367), .B(n1863), .CI(n1356), .CO(n1349), .S(n1350) );
  ADD32 U729 ( .A(n1803), .B(n1893), .CI(n1833), .CO(n1351), .S(n1352) );
  ADD32 U730 ( .A(n1743), .B(n1923), .CI(n1773), .CO(n1353), .S(n1354) );
  ADD22 U731 ( .A(n1449), .B(n1954), .CO(n1355), .S(n1356) );
  ADD32 U732 ( .A(n1371), .B(n1362), .CI(n1360), .CO(n1357), .S(n1358) );
  ADD32 U733 ( .A(n1373), .B(n1366), .CI(n1364), .CO(n1359), .S(n1360) );
  ADD32 U734 ( .A(n1375), .B(n1377), .CI(n1368), .CO(n1361), .S(n1362) );
  ADD32 U735 ( .A(n1834), .B(n1864), .CI(n1379), .CO(n1363), .S(n1364) );
  ADD32 U736 ( .A(n1804), .B(n1894), .CI(n1744), .CO(n1365), .S(n1366) );
  ADD32 U737 ( .A(n1924), .B(n1955), .CI(n1774), .CO(n1367), .S(n1368) );
  ADD32 U738 ( .A(n1383), .B(n1374), .CI(n1372), .CO(n1369), .S(n1370) );
  ADD32 U739 ( .A(n1378), .B(n1376), .CI(n1385), .CO(n1371), .S(n1372) );
  ADD32 U740 ( .A(n1380), .B(n1389), .CI(n1387), .CO(n1373), .S(n1374) );
  ADD32 U741 ( .A(n1805), .B(n1865), .CI(n1835), .CO(n1375), .S(n1376) );
  ADD32 U742 ( .A(n1775), .B(n1925), .CI(n1895), .CO(n1377), .S(n1378) );
  ADD22 U743 ( .A(n1450), .B(n1956), .CO(n1379), .S(n1380) );
  ADD32 U744 ( .A(n1393), .B(n1386), .CI(n1384), .CO(n1381), .S(n1382) );
  ADD32 U745 ( .A(n1388), .B(n1390), .CI(n1395), .CO(n1383), .S(n1384) );
  ADD32 U746 ( .A(n1399), .B(n1866), .CI(n1397), .CO(n1385), .S(n1386) );
  ADD32 U747 ( .A(n1836), .B(n1896), .CI(n1776), .CO(n1387), .S(n1388) );
  ADD32 U748 ( .A(n1926), .B(n1957), .CI(n1806), .CO(n1389), .S(n1390) );
  ADD32 U749 ( .A(n1403), .B(n1396), .CI(n1394), .CO(n1391), .S(n1392) );
  ADD32 U750 ( .A(n1405), .B(n1400), .CI(n1398), .CO(n1393), .S(n1394) );
  ADD32 U751 ( .A(n1837), .B(n1867), .CI(n1407), .CO(n1395), .S(n1396) );
  ADD32 U752 ( .A(n1807), .B(n1927), .CI(n1897), .CO(n1397), .S(n1398) );
  ADD22 U753 ( .A(n1451), .B(n1958), .CO(n1399), .S(n1400) );
  ADD32 U754 ( .A(n1411), .B(n1406), .CI(n1404), .CO(n1401), .S(n1402) );
  ADD32 U755 ( .A(n1413), .B(n1415), .CI(n1408), .CO(n1403), .S(n1404) );
  ADD32 U756 ( .A(n1868), .B(n1898), .CI(n1808), .CO(n1405), .S(n1406) );
  ADD32 U757 ( .A(n1928), .B(n1959), .CI(n1838), .CO(n1407), .S(n1408) );
  ADD32 U758 ( .A(n1419), .B(n1414), .CI(n1412), .CO(n1409), .S(n1410) );
  ADD32 U759 ( .A(n1421), .B(n1899), .CI(n1416), .CO(n1411), .S(n1412) );
  ADD32 U760 ( .A(n1839), .B(n1929), .CI(n1869), .CO(n1413), .S(n1414) );
  ADD22 U761 ( .A(n1452), .B(n1960), .CO(n1415), .S(n1416) );
  ADD32 U762 ( .A(n1422), .B(n1425), .CI(n1420), .CO(n1417), .S(n1418) );
  ADD32 U763 ( .A(n1840), .B(n1900), .CI(n1427), .CO(n1419), .S(n1420) );
  ADD32 U764 ( .A(n1930), .B(n1961), .CI(n1870), .CO(n1421), .S(n1422) );
  ADD32 U765 ( .A(n1428), .B(n1431), .CI(n1426), .CO(n1423), .S(n1424) );
  ADD32 U766 ( .A(n1871), .B(n1931), .CI(n1901), .CO(n1425), .S(n1426) );
  ADD22 U767 ( .A(n1453), .B(n1962), .CO(n1427), .S(n1428) );
  ADD32 U768 ( .A(n1435), .B(n1872), .CI(n1432), .CO(n1429), .S(n1430) );
  ADD32 U769 ( .A(n1932), .B(n1963), .CI(n1902), .CO(n1431), .S(n1432) );
  ADD32 U770 ( .A(n1903), .B(n1933), .CI(n1437), .CO(n1433), .S(n1434) );
  ADD22 U771 ( .A(n1454), .B(n1964), .CO(n1435), .S(n1436) );
  ADD32 U772 ( .A(n1934), .B(n1965), .CI(n1904), .CO(n1437), .S(n1438) );
  ADD22 U773 ( .A(n1935), .B(n1966), .CO(n1439), .S(n1440) );
  OAI222 U1910 ( .A(n3060), .B(n2997), .C(n2816), .D(n3061), .Q(n1932) );
  CLKBU12 U1911 ( .A(n2980), .Q(n2815) );
  INV12 U1912 ( .A(a[0]), .Q(n2985) );
  XNR21 U1913 ( .A(n2818), .B(n2892), .Q(n3025) );
  NAND33 U1914 ( .A(n2750), .B(n2751), .C(n2752), .Q(n504) );
  NAND33 U1915 ( .A(n2783), .B(n2784), .C(n2785), .Q(n469) );
  NAND33 U1916 ( .A(n2780), .B(n2781), .C(n2782), .Q(n459) );
  CLKIN8 U1917 ( .A(a[3]), .Q(n2897) );
  NAND32 U1918 ( .A(n2810), .B(n2811), .C(n2812), .Q(n450) );
  NAND22 U1919 ( .A(n3522), .B(n2986), .Q(n3521) );
  OAI221 U1920 ( .A(n2940), .B(n3508), .C(n3507), .D(n3023), .Q(n1467) );
  AOI211 U1921 ( .A(n2999), .B(n3521), .C(n2900), .Q(n1454) );
  OAI221 U1922 ( .A(n2940), .B(n3510), .C(n3509), .D(n3023), .Q(n1465) );
  OAI221 U1923 ( .A(n2980), .B(n3089), .C(n3088), .D(n2999), .Q(n1903) );
  OAI221 U1924 ( .A(n2940), .B(n3511), .C(n3510), .D(n3023), .Q(n1464) );
  NAND22 U1925 ( .A(n2959), .B(n3544), .Q(n3012) );
  OAI221 U1926 ( .A(n2962), .B(n2742), .C(n3009), .D(n3010), .Q(n637) );
  OAI221 U1927 ( .A(n2940), .B(n3512), .C(n3511), .D(n3023), .Q(n1463) );
  XNR21 U1928 ( .A(n2986), .B(n2900), .Q(n3088) );
  NAND22 U1929 ( .A(n2968), .B(n3535), .Q(n2994) );
  OAI221 U1930 ( .A(n2953), .B(n2745), .C(n3015), .D(n3016), .Q(n559) );
  OAI221 U1931 ( .A(n2940), .B(n3513), .C(n3512), .D(n3023), .Q(n1462) );
  NAND22 U1932 ( .A(n2971), .B(n3532), .Q(n3005) );
  OAI221 U1933 ( .A(n2968), .B(n3214), .C(n3213), .D(n2994), .Q(n1774) );
  OAI221 U1934 ( .A(n2940), .B(n3509), .C(n3508), .D(n3023), .Q(n1466) );
  OAI221 U1935 ( .A(n2944), .B(n2748), .C(n3021), .D(n2991), .Q(n517) );
  NOR22 U1936 ( .A(n2977), .B(n2986), .Q(n1872) );
  NAND34 U1937 ( .A(n2773), .B(n2774), .C(n2775), .Q(n503) );
  NAND34 U1938 ( .A(n2792), .B(n2793), .C(n2794), .Q(n502) );
  XNR21 U1939 ( .A(a[4]), .B(n2897), .Q(n3522) );
  NAND32 U1940 ( .A(n2758), .B(n2759), .C(n2760), .Q(n508) );
  NAND33 U1941 ( .A(n2807), .B(n2808), .C(n2809), .Q(n501) );
  NAND22 U1942 ( .A(n1402), .B(n1409), .Q(n2809) );
  XOR21 U1943 ( .A(n450), .B(n2776), .Q(product[62]) );
  INV6 U1944 ( .A(n3519), .Q(n2983) );
  NAND24 U1945 ( .A(n459), .B(n561), .Q(n2796) );
  NAND24 U1946 ( .A(n459), .B(n552), .Q(n2795) );
  OAI222 U1947 ( .A(n3091), .B(n2859), .C(n2814), .D(n3092), .Q(n1900) );
  OAI222 U1948 ( .A(b[0]), .B(n3024), .C(n3025), .D(n2985), .Q(n1968) );
  OAI222 U1949 ( .A(n3025), .B(n2756), .C(n3026), .D(n2985), .Q(n1967) );
  XOR21 U1950 ( .A(a[6]), .B(a[5]), .Q(n3525) );
  BUF6 U1951 ( .A(n2983), .Q(n2816) );
  CLKIN6 U1952 ( .A(n2894), .Q(n2892) );
  CLKBU6 U1953 ( .A(n2983), .Q(n2817) );
  NAND32 U1954 ( .A(n2789), .B(n2790), .C(n2791), .Q(n489) );
  NAND32 U1955 ( .A(n2786), .B(n2787), .C(n2788), .Q(n479) );
  NAND22 U1956 ( .A(n2892), .B(n2985), .Q(n3024) );
  NAND22 U1957 ( .A(n2815), .B(n3523), .Q(n2999) );
  NAND22 U1958 ( .A(n2817), .B(n3520), .Q(n2997) );
  XOR21 U1959 ( .A(n2848), .B(n2908), .Q(n2739) );
  XOR21 U1960 ( .A(n2848), .B(n2910), .Q(n2740) );
  XOR21 U1961 ( .A(n2848), .B(n2913), .Q(n2741) );
  XOR21 U1962 ( .A(n2848), .B(n2916), .Q(n2742) );
  XOR21 U1963 ( .A(n2848), .B(n2919), .Q(n2743) );
  XOR21 U1964 ( .A(n2848), .B(n2922), .Q(n2744) );
  XOR21 U1965 ( .A(n2848), .B(n2924), .Q(n2745) );
  XOR21 U1966 ( .A(n2848), .B(n2927), .Q(n2746) );
  XOR21 U1967 ( .A(n2848), .B(n2930), .Q(n2747) );
  XOR21 U1968 ( .A(n2848), .B(n2933), .Q(n2748) );
  XOR21 U1969 ( .A(n2848), .B(n2936), .Q(n2749) );
  CLKIN6 U1970 ( .A(a[1]), .Q(n2894) );
  XOR21 U1971 ( .A(a[8]), .B(a[7]), .Q(n3528) );
  NAND24 U1972 ( .A(n469), .B(n711), .Q(n2799) );
  XOR31 U1973 ( .A(n505), .B(n1424), .C(n1429), .Q(product[7]) );
  NAND22 U1974 ( .A(n505), .B(n1424), .Q(n2750) );
  NAND22 U1975 ( .A(n505), .B(n1429), .Q(n2751) );
  NAND22 U1976 ( .A(n1424), .B(n1429), .Q(n2752) );
  NAND33 U1977 ( .A(n2767), .B(n2768), .C(n2769), .Q(n480) );
  NAND33 U1978 ( .A(n2764), .B(n2765), .C(n2766), .Q(n470) );
  NAND33 U1979 ( .A(n2770), .B(n2771), .C(n2772), .Q(n490) );
  NAND33 U1980 ( .A(n2761), .B(n2762), .C(n2763), .Q(n460) );
  NAND33 U1981 ( .A(n2798), .B(n2799), .C(n2800), .Q(n468) );
  XOR21 U1982 ( .A(n2848), .B(n2900), .Q(n2753) );
  XOR21 U1983 ( .A(n2848), .B(n2903), .Q(n2754) );
  XOR21 U1984 ( .A(n2848), .B(n2906), .Q(n2755) );
  NAND22 U1985 ( .A(n2892), .B(n2985), .Q(n2756) );
  NAND22 U1986 ( .A(n992), .B(n1021), .Q(n2769) );
  NAND22 U1987 ( .A(n481), .B(n1021), .Q(n2768) );
  NAND22 U1988 ( .A(n481), .B(n992), .Q(n2767) );
  NAND22 U1989 ( .A(n732), .B(n753), .Q(n2766) );
  NAND22 U1990 ( .A(n471), .B(n753), .Q(n2765) );
  NAND22 U1991 ( .A(n471), .B(n732), .Q(n2764) );
  NAND22 U1992 ( .A(n731), .B(n712), .Q(n2785) );
  NAND22 U1993 ( .A(n470), .B(n712), .Q(n2784) );
  NAND22 U1994 ( .A(n470), .B(n731), .Q(n2783) );
  NAND22 U1995 ( .A(n1242), .B(n1261), .Q(n2772) );
  NAND22 U1996 ( .A(n491), .B(n1261), .Q(n2771) );
  NAND22 U1997 ( .A(n491), .B(n1242), .Q(n2770) );
  NAND22 U1998 ( .A(n1222), .B(n1241), .Q(n2791) );
  NAND22 U1999 ( .A(n490), .B(n1241), .Q(n2790) );
  NAND22 U2000 ( .A(n490), .B(n1222), .Q(n2789) );
  NAND22 U2001 ( .A(n962), .B(n991), .Q(n2788) );
  NAND22 U2002 ( .A(n480), .B(n991), .Q(n2787) );
  NAND22 U2003 ( .A(n480), .B(n962), .Q(n2786) );
  NAND22 U2004 ( .A(n572), .B(n583), .Q(n2763) );
  NAND22 U2005 ( .A(n461), .B(n583), .Q(n2762) );
  NAND22 U2006 ( .A(n461), .B(n572), .Q(n2761) );
  NAND33 U2007 ( .A(n2804), .B(n2805), .C(n2806), .Q(n488) );
  NAND22 U2008 ( .A(n1200), .B(n1221), .Q(n2806) );
  NAND22 U2009 ( .A(n489), .B(n1200), .Q(n2804) );
  NAND33 U2010 ( .A(n2801), .B(n2802), .C(n2803), .Q(n478) );
  NAND22 U2011 ( .A(n932), .B(n961), .Q(n2803) );
  NAND22 U2012 ( .A(n479), .B(n932), .Q(n2801) );
  NAND22 U2013 ( .A(n692), .B(n711), .Q(n2800) );
  NAND22 U2014 ( .A(n489), .B(n1221), .Q(n2805) );
  NAND22 U2015 ( .A(n479), .B(n961), .Q(n2802) );
  NAND22 U2016 ( .A(n571), .B(n562), .Q(n2782) );
  NAND22 U2017 ( .A(n460), .B(n562), .Q(n2781) );
  NAND22 U2018 ( .A(n460), .B(n571), .Q(n2780) );
  NAND33 U2019 ( .A(n2795), .B(n2796), .C(n2797), .Q(n458) );
  NAND22 U2020 ( .A(n552), .B(n561), .Q(n2797) );
  NAND22 U2021 ( .A(n1418), .B(n1423), .Q(n2775) );
  NAND22 U2022 ( .A(n1410), .B(n1417), .Q(n2794) );
  NAND32 U2023 ( .A(n2777), .B(n2778), .C(n2779), .Q(n449) );
  CLKIN6 U2024 ( .A(n511), .Q(n2938) );
  CLKBU6 U2025 ( .A(n2980), .Q(n2814) );
  CLKBU6 U2026 ( .A(n2977), .Q(n2813) );
  CLKBU6 U2027 ( .A(n2756), .Q(n2891) );
  OAI221 U2028 ( .A(n3022), .B(n3023), .C(n2940), .D(n2749), .Q(n511) );
  OAI221 U2029 ( .A(n3057), .B(n2997), .C(n2817), .D(n3058), .Q(n1935) );
  CLKIN6 U2030 ( .A(n3522), .Q(n2980) );
  CLKIN6 U2031 ( .A(n3525), .Q(n2977) );
  CLKIN6 U2032 ( .A(n3531), .Q(n2971) );
  CLKIN6 U2033 ( .A(n3528), .Q(n2974) );
  CLKIN6 U2034 ( .A(n2897), .Q(n2895) );
  CLKIN6 U2035 ( .A(n2894), .Q(n2893) );
  CLKIN6 U2036 ( .A(n2903), .Q(n2901) );
  CLKIN6 U2037 ( .A(n2900), .Q(n2898) );
  CLKBU6 U2038 ( .A(n2997), .Q(n2857) );
  CLKIN6 U2039 ( .A(n3534), .Q(n2968) );
  CLKIN6 U2040 ( .A(n3537), .Q(n2965) );
  CLKIN6 U2041 ( .A(n2906), .Q(n2904) );
  CLKIN6 U2042 ( .A(n2908), .Q(n2907) );
  CLKBU6 U2043 ( .A(n3001), .Q(n2861) );
  CLKIN6 U2044 ( .A(n2897), .Q(n2896) );
  CLKIN6 U2045 ( .A(n2910), .Q(n2909) );
  CLKBU6 U2046 ( .A(n3003), .Q(n2862) );
  CLKIN6 U2047 ( .A(n3540), .Q(n2962) );
  CLKIN6 U2048 ( .A(n2900), .Q(n2899) );
  CLKBU6 U2049 ( .A(n3010), .Q(n2865) );
  CLKBU6 U2050 ( .A(n3005), .Q(n2863) );
  CLKBU6 U2051 ( .A(n2994), .Q(n2856) );
  CLKBU6 U2052 ( .A(n2997), .Q(n2858) );
  CLKBU6 U2053 ( .A(n2986), .Q(n2849) );
  CLKIN6 U2054 ( .A(n3543), .Q(n2959) );
  CLKIN6 U2055 ( .A(n2903), .Q(n2902) );
  CLKIN6 U2056 ( .A(n2913), .Q(n2911) );
  CLKIN6 U2057 ( .A(n2916), .Q(n2914) );
  CLKBU6 U2058 ( .A(n2999), .Q(n2859) );
  CLKIN6 U2059 ( .A(n3549), .Q(n2953) );
  CLKIN6 U2060 ( .A(n3546), .Q(n2956) );
  CLKIN6 U2061 ( .A(n2906), .Q(n2905) );
  CLKBU6 U2062 ( .A(n2986), .Q(n2850) );
  CLKBU6 U2063 ( .A(n3016), .Q(n2876) );
  CLKBU6 U2064 ( .A(n3014), .Q(n2871) );
  CLKIN6 U2065 ( .A(n2919), .Q(n2917) );
  CLKIN6 U2066 ( .A(n2922), .Q(n2920) );
  CLKBU6 U2067 ( .A(n3010), .Q(n2866) );
  CLKBU6 U2068 ( .A(n2999), .Q(n2860) );
  CLKIN6 U2069 ( .A(n3552), .Q(n2950) );
  CLKIN6 U2070 ( .A(n3555), .Q(n2947) );
  CLKIN6 U2071 ( .A(n2924), .Q(n2923) );
  CLKBU6 U2072 ( .A(n3018), .Q(n2881) );
  CLKIN6 U2073 ( .A(n3558), .Q(n2944) );
  CLKIN6 U2074 ( .A(n2913), .Q(n2912) );
  CLKIN6 U2075 ( .A(n2927), .Q(n2925) );
  CLKBU6 U2076 ( .A(n3014), .Q(n2872) );
  CLKBU6 U2077 ( .A(n2991), .Q(n2851) );
  CLKIN6 U2078 ( .A(n3561), .Q(n2940) );
  CLKIN6 U2079 ( .A(n2916), .Q(n2915) );
  CLKIN6 U2080 ( .A(n2930), .Q(n2928) );
  CLKBU6 U2081 ( .A(n3016), .Q(n2877) );
  CLKBU6 U2082 ( .A(n3010), .Q(n2867) );
  CLKIN6 U2083 ( .A(n2919), .Q(n2918) );
  CLKBU6 U2084 ( .A(n3018), .Q(n2882) );
  CLKBU6 U2085 ( .A(n3020), .Q(n2886) );
  CLKIN6 U2086 ( .A(n2922), .Q(n2921) );
  CLKIN6 U2087 ( .A(n2933), .Q(n2931) );
  CLKIN6 U2088 ( .A(n2936), .Q(n2934) );
  CLKBU6 U2089 ( .A(n2991), .Q(n2853) );
  XOR21 U2090 ( .A(n2848), .B(n2897), .Q(n2757) );
  CLKBU6 U2091 ( .A(n3016), .Q(n2878) );
  CLKBU6 U2092 ( .A(n3014), .Q(n2873) );
  CLKBU6 U2093 ( .A(n2991), .Q(n2852) );
  CLKIN6 U2094 ( .A(n2927), .Q(n2926) );
  CLKBU6 U2095 ( .A(n3010), .Q(n2868) );
  CLKIN6 U2096 ( .A(n2930), .Q(n2929) );
  CLKBU6 U2097 ( .A(n3018), .Q(n2883) );
  CLKIN6 U2098 ( .A(n2933), .Q(n2932) );
  CLKBU6 U2099 ( .A(n3020), .Q(n2887) );
  CLKBU6 U2100 ( .A(n3014), .Q(n2874) );
  CLKBU6 U2101 ( .A(n3008), .Q(n2864) );
  CLKIN6 U2102 ( .A(n2936), .Q(n2935) );
  CLKBU6 U2103 ( .A(n3016), .Q(n2879) );
  CLKBU6 U2104 ( .A(n3010), .Q(n2869) );
  CLKBU6 U2105 ( .A(n3018), .Q(n2884) );
  CLKBU6 U2106 ( .A(n3012), .Q(n2870) );
  CLKBU6 U2107 ( .A(n3020), .Q(n2888) );
  CLKBU6 U2108 ( .A(n3014), .Q(n2875) );
  CLKBU6 U2109 ( .A(n2991), .Q(n2854) );
  CLKBU6 U2110 ( .A(n3016), .Q(n2880) );
  CLKBU6 U2111 ( .A(n3018), .Q(n2885) );
  CLKBU6 U2112 ( .A(n2991), .Q(n2855) );
  CLKBU6 U2113 ( .A(n3020), .Q(n2889) );
  CLKBU6 U2114 ( .A(n3023), .Q(n2890) );
  NAND22 U2115 ( .A(n2977), .B(n3526), .Q(n3001) );
  CLKBU6 U2116 ( .A(b[6]), .Q(n2823) );
  CLKBU6 U2117 ( .A(b[3]), .Q(n2820) );
  CLKBU6 U2118 ( .A(b[4]), .Q(n2821) );
  CLKBU6 U2119 ( .A(b[2]), .Q(n2819) );
  CLKBU6 U2120 ( .A(b[1]), .Q(n2818) );
  XNR21 U2121 ( .A(a[2]), .B(n2897), .Q(n3520) );
  CLKIN6 U2122 ( .A(a[9]), .Q(n2906) );
  CLKIN6 U2123 ( .A(a[7]), .Q(n2903) );
  CLKIN6 U2124 ( .A(a[5]), .Q(n2900) );
  CLKBU6 U2125 ( .A(b[5]), .Q(n2822) );
  CLKBU6 U2126 ( .A(b[7]), .Q(n2824) );
  CLKIN6 U2127 ( .A(a[11]), .Q(n2908) );
  CLKBU6 U2128 ( .A(b[8]), .Q(n2825) );
  CLKBU6 U2129 ( .A(b[9]), .Q(n2826) );
  CLKBU6 U2130 ( .A(b[10]), .Q(n2827) );
  CLKBU6 U2131 ( .A(b[11]), .Q(n2828) );
  CLKIN6 U2132 ( .A(a[13]), .Q(n2910) );
  CLKBU6 U2133 ( .A(b[12]), .Q(n2829) );
  CLKIN6 U2134 ( .A(a[15]), .Q(n2913) );
  CLKBU6 U2135 ( .A(b[15]), .Q(n2832) );
  CLKBU6 U2136 ( .A(b[13]), .Q(n2830) );
  CLKBU6 U2137 ( .A(b[14]), .Q(n2831) );
  CLKBU6 U2138 ( .A(b[16]), .Q(n2833) );
  CLKBU6 U2139 ( .A(b[17]), .Q(n2834) );
  CLKBU6 U2140 ( .A(b[18]), .Q(n2835) );
  CLKIN6 U2141 ( .A(a[17]), .Q(n2916) );
  CLKBU6 U2142 ( .A(b[19]), .Q(n2836) );
  CLKIN6 U2143 ( .A(a[19]), .Q(n2919) );
  CLKIN6 U2144 ( .A(a[21]), .Q(n2922) );
  CLKBU6 U2145 ( .A(b[20]), .Q(n2837) );
  CLKIN6 U2146 ( .A(a[23]), .Q(n2924) );
  CLKBU6 U2147 ( .A(b[21]), .Q(n2838) );
  CLKBU6 U2148 ( .A(b[22]), .Q(n2839) );
  CLKBU6 U2149 ( .A(b[23]), .Q(n2840) );
  CLKIN6 U2150 ( .A(a[25]), .Q(n2927) );
  CLKBU6 U2151 ( .A(b[24]), .Q(n2841) );
  CLKIN6 U2152 ( .A(a[27]), .Q(n2930) );
  CLKBU6 U2153 ( .A(b[28]), .Q(n2845) );
  CLKBU6 U2154 ( .A(b[27]), .Q(n2844) );
  CLKBU6 U2155 ( .A(b[25]), .Q(n2842) );
  CLKBU6 U2156 ( .A(b[26]), .Q(n2843) );
  CLKIN6 U2157 ( .A(a[29]), .Q(n2933) );
  CLKBU6 U2158 ( .A(b[29]), .Q(n2846) );
  CLKBU6 U2159 ( .A(b[30]), .Q(n2847) );
  CLKBU6 U2160 ( .A(b[31]), .Q(n2848) );
  CLKIN6 U2161 ( .A(a[31]), .Q(n2936) );
  XOR31 U2162 ( .A(n1440), .B(n509), .C(n1455), .Q(product[3]) );
  NAND22 U2163 ( .A(n509), .B(n1440), .Q(n2758) );
  NAND22 U2164 ( .A(n1440), .B(n1455), .Q(n2759) );
  NAND22 U2165 ( .A(n509), .B(n1455), .Q(n2760) );
  XOR31 U2166 ( .A(n461), .B(n572), .C(n583), .Q(product[51]) );
  XOR31 U2167 ( .A(n471), .B(n732), .C(n753), .Q(product[41]) );
  XOR31 U2168 ( .A(n481), .B(n992), .C(n1021), .Q(product[31]) );
  XOR31 U2169 ( .A(n491), .B(n1242), .C(n1261), .Q(product[21]) );
  XOR31 U2170 ( .A(n504), .B(n1418), .C(n1423), .Q(product[8]) );
  NAND24 U2171 ( .A(n504), .B(n1418), .Q(n2773) );
  NAND24 U2172 ( .A(n504), .B(n1423), .Q(n2774) );
  XOR21 U2173 ( .A(n511), .B(n2939), .Q(n2776) );
  NAND22 U2174 ( .A(n450), .B(n511), .Q(n2777) );
  NAND22 U2175 ( .A(n450), .B(n2939), .Q(n2778) );
  NAND22 U2176 ( .A(n511), .B(n2939), .Q(n2779) );
  XOR31 U2177 ( .A(n460), .B(n571), .C(n562), .Q(product[52]) );
  XOR31 U2178 ( .A(n470), .B(n731), .C(n712), .Q(product[42]) );
  XOR31 U2179 ( .A(n480), .B(n962), .C(n991), .Q(product[32]) );
  XOR31 U2180 ( .A(n490), .B(n1222), .C(n1241), .Q(product[22]) );
  XOR31 U2181 ( .A(n503), .B(n1410), .C(n1417), .Q(product[9]) );
  NAND24 U2182 ( .A(n503), .B(n1410), .Q(n2792) );
  NAND24 U2183 ( .A(n503), .B(n1417), .Q(n2793) );
  OAI222 U2184 ( .A(n3089), .B(n2999), .C(n2814), .D(n3090), .Q(n1902) );
  XNR22 U2185 ( .A(a[2]), .B(n2894), .Q(n3519) );
  XOR31 U2186 ( .A(n459), .B(n552), .C(n561), .Q(product[53]) );
  XOR31 U2187 ( .A(n469), .B(n692), .C(n711), .Q(product[43]) );
  NAND24 U2188 ( .A(n469), .B(n692), .Q(n2798) );
  XOR31 U2189 ( .A(n479), .B(n932), .C(n961), .Q(product[33]) );
  XOR31 U2190 ( .A(n489), .B(n1200), .C(n1221), .Q(product[23]) );
  XOR31 U2191 ( .A(n502), .B(n1402), .C(n1409), .Q(product[10]) );
  NAND24 U2192 ( .A(n502), .B(n1402), .Q(n2807) );
  NAND24 U2193 ( .A(n502), .B(n1409), .Q(n2808) );
  XOR31 U2194 ( .A(n451), .B(n513), .C(n2938), .Q(product[61]) );
  NAND22 U2195 ( .A(n451), .B(n513), .Q(n2810) );
  NAND22 U2196 ( .A(n451), .B(n2938), .Q(n2811) );
  NAND22 U2197 ( .A(n513), .B(n2938), .Q(n2812) );
  CLKIN6 U2198 ( .A(n449), .Q(product[63]) );
  CLKIN6 U2199 ( .A(n3517), .Q(n2939) );
  CLKIN6 U2200 ( .A(n2989), .Q(n2941) );
  CLKIN6 U2201 ( .A(n517), .Q(n2942) );
  CLKIN6 U2202 ( .A(n3486), .Q(n2943) );
  CLKIN6 U2203 ( .A(n527), .Q(n2945) );
  CLKIN6 U2204 ( .A(n3457), .Q(n2946) );
  CLKIN6 U2205 ( .A(n541), .Q(n2948) );
  CLKIN6 U2206 ( .A(n3426), .Q(n2949) );
  CLKIN6 U2207 ( .A(n559), .Q(n2951) );
  CLKIN6 U2208 ( .A(n3395), .Q(n2952) );
  CLKIN6 U2209 ( .A(n581), .Q(n2954) );
  CLKIN6 U2210 ( .A(n3364), .Q(n2955) );
  CLKIN6 U2211 ( .A(n607), .Q(n2957) );
  CLKIN6 U2212 ( .A(n3333), .Q(n2958) );
  CLKIN6 U2213 ( .A(n637), .Q(n2960) );
  CLKIN6 U2214 ( .A(n3302), .Q(n2961) );
  CLKIN6 U2215 ( .A(n671), .Q(n2963) );
  CLKIN6 U2216 ( .A(n3271), .Q(n2964) );
  CLKIN6 U2217 ( .A(n709), .Q(n2966) );
  CLKIN6 U2218 ( .A(n3240), .Q(n2967) );
  CLKIN6 U2219 ( .A(n751), .Q(n2969) );
  CLKIN6 U2220 ( .A(n3211), .Q(n2970) );
  CLKIN6 U2221 ( .A(n797), .Q(n2972) );
  CLKIN6 U2222 ( .A(n3180), .Q(n2973) );
  CLKIN6 U2223 ( .A(n847), .Q(n2975) );
  CLKIN6 U2224 ( .A(n3149), .Q(n2976) );
  CLKIN6 U2225 ( .A(n901), .Q(n2978) );
  CLKIN6 U2226 ( .A(n3118), .Q(n2979) );
  CLKIN6 U2227 ( .A(n959), .Q(n2981) );
  CLKIN6 U2228 ( .A(n3087), .Q(n2982) );
  CLKIN6 U2229 ( .A(n3056), .Q(n2984) );
  CLKIN6 U2230 ( .A(b[0]), .Q(n2986) );
  NOR22 U2231 ( .A(n2849), .B(n2985), .Q(product[0]) );
  XNR21 U2232 ( .A(n2987), .B(n2988), .Q(n990) );
  NOR22 U2233 ( .A(n2988), .B(n2987), .Q(n2989) );
  OAI221 U2234 ( .A(n2990), .B(n2853), .C(n2944), .D(n2992), .Q(n2987) );
  OAI221 U2235 ( .A(n2993), .B(n2856), .C(n2968), .D(n2995), .Q(n2988) );
  OAI221 U2236 ( .A(n2996), .B(n2858), .C(n2816), .D(n2757), .Q(n959) );
  OAI221 U2237 ( .A(n2998), .B(n2859), .C(n2814), .D(n2753), .Q(n901) );
  OAI221 U2238 ( .A(n3000), .B(n2861), .C(n2813), .D(n2754), .Q(n847) );
  OAI221 U2239 ( .A(n3002), .B(n2862), .C(n2974), .D(n2755), .Q(n797) );
  OAI221 U2240 ( .A(n3004), .B(n2863), .C(n2971), .D(n2739), .Q(n751) );
  OAI221 U2241 ( .A(n3006), .B(n2856), .C(n2968), .D(n2740), .Q(n709) );
  OAI221 U2242 ( .A(n3007), .B(n2864), .C(n2965), .D(n2741), .Q(n671) );
  OAI221 U2243 ( .A(n3011), .B(n2870), .C(n2959), .D(n2743), .Q(n607) );
  OAI221 U2244 ( .A(n3013), .B(n2873), .C(n2956), .D(n2744), .Q(n581) );
  OAI221 U2245 ( .A(n3017), .B(n2883), .C(n2950), .D(n2746), .Q(n541) );
  OAI221 U2246 ( .A(n3019), .B(n2887), .C(n2947), .D(n2747), .Q(n527) );
  OAI221 U2247 ( .A(n3026), .B(n2756), .C(n3027), .D(n2985), .Q(n1966) );
  XNR21 U2248 ( .A(n2819), .B(n2892), .Q(n3026) );
  OAI221 U2249 ( .A(n3027), .B(n2756), .C(n3028), .D(n2985), .Q(n1965) );
  XNR21 U2250 ( .A(n2820), .B(n2892), .Q(n3027) );
  OAI221 U2251 ( .A(n3028), .B(n2891), .C(n3029), .D(n2985), .Q(n1964) );
  XNR21 U2252 ( .A(n2821), .B(n2892), .Q(n3028) );
  OAI221 U2253 ( .A(n3029), .B(n2756), .C(n3030), .D(n2985), .Q(n1963) );
  XNR21 U2254 ( .A(n2822), .B(n2892), .Q(n3029) );
  OAI221 U2255 ( .A(n3030), .B(n2891), .C(n3031), .D(n2985), .Q(n1962) );
  XNR21 U2256 ( .A(n2823), .B(n2892), .Q(n3030) );
  OAI221 U2257 ( .A(n3031), .B(n2756), .C(n3032), .D(n2985), .Q(n1961) );
  XNR21 U2258 ( .A(n2824), .B(n2892), .Q(n3031) );
  OAI221 U2259 ( .A(n3032), .B(n2756), .C(n3033), .D(n2985), .Q(n1960) );
  XNR21 U2260 ( .A(n2825), .B(n2892), .Q(n3032) );
  OAI221 U2261 ( .A(n3033), .B(n2891), .C(n3034), .D(n2985), .Q(n1959) );
  XNR21 U2262 ( .A(n2826), .B(n2892), .Q(n3033) );
  OAI221 U2263 ( .A(n3034), .B(n2891), .C(n3035), .D(n2985), .Q(n1958) );
  XNR21 U2264 ( .A(n2827), .B(n2893), .Q(n3034) );
  OAI221 U2265 ( .A(n3035), .B(n2891), .C(n3036), .D(n2985), .Q(n1957) );
  XNR21 U2266 ( .A(n2828), .B(n2893), .Q(n3035) );
  OAI221 U2267 ( .A(n3036), .B(n2891), .C(n3037), .D(n2985), .Q(n1956) );
  XNR21 U2268 ( .A(n2829), .B(n2893), .Q(n3036) );
  OAI221 U2269 ( .A(n3037), .B(n2891), .C(n3038), .D(n2985), .Q(n1955) );
  XNR21 U2270 ( .A(n2830), .B(n2893), .Q(n3037) );
  OAI221 U2271 ( .A(n3038), .B(n2891), .C(n3039), .D(n2985), .Q(n1954) );
  XNR21 U2272 ( .A(n2831), .B(n2893), .Q(n3038) );
  OAI221 U2273 ( .A(n3039), .B(n2891), .C(n3040), .D(n2985), .Q(n1953) );
  XNR21 U2274 ( .A(n2832), .B(n2893), .Q(n3039) );
  OAI221 U2275 ( .A(n3040), .B(n2891), .C(n3041), .D(n2985), .Q(n1952) );
  XNR21 U2276 ( .A(n2833), .B(n2893), .Q(n3040) );
  OAI221 U2277 ( .A(n3041), .B(n2891), .C(n3042), .D(n2985), .Q(n1951) );
  XNR21 U2278 ( .A(n2834), .B(n2893), .Q(n3041) );
  OAI221 U2279 ( .A(n3042), .B(n2891), .C(n3043), .D(n2985), .Q(n1950) );
  XNR21 U2280 ( .A(n2835), .B(n2893), .Q(n3042) );
  OAI221 U2281 ( .A(n3043), .B(n2891), .C(n3044), .D(n2985), .Q(n1949) );
  XNR21 U2282 ( .A(n2836), .B(n2893), .Q(n3043) );
  OAI221 U2283 ( .A(n3044), .B(n2891), .C(n3045), .D(n2985), .Q(n1948) );
  XNR21 U2284 ( .A(n2837), .B(n2893), .Q(n3044) );
  OAI221 U2285 ( .A(n3045), .B(n2891), .C(n3046), .D(n2985), .Q(n1947) );
  XNR21 U2286 ( .A(n2838), .B(n2893), .Q(n3045) );
  OAI221 U2287 ( .A(n3046), .B(n2891), .C(n3047), .D(n2985), .Q(n1946) );
  XNR21 U2288 ( .A(n2839), .B(n2893), .Q(n3046) );
  OAI221 U2289 ( .A(n3047), .B(n2891), .C(n3048), .D(n2985), .Q(n1945) );
  XNR21 U2290 ( .A(n2840), .B(n2893), .Q(n3047) );
  OAI221 U2291 ( .A(n3048), .B(n2891), .C(n3049), .D(n2985), .Q(n1944) );
  XNR21 U2292 ( .A(n2841), .B(n2893), .Q(n3048) );
  OAI221 U2293 ( .A(n3049), .B(n2891), .C(n3050), .D(n2985), .Q(n1943) );
  XNR21 U2294 ( .A(n2842), .B(n2893), .Q(n3049) );
  OAI221 U2295 ( .A(n3050), .B(n2891), .C(n3051), .D(n2985), .Q(n1942) );
  XNR21 U2296 ( .A(n2843), .B(n2893), .Q(n3050) );
  OAI221 U2297 ( .A(n3051), .B(n2891), .C(n3052), .D(n2985), .Q(n1941) );
  XNR21 U2298 ( .A(n2844), .B(n2893), .Q(n3051) );
  OAI221 U2299 ( .A(n3052), .B(n2891), .C(n3053), .D(n2985), .Q(n1940) );
  XNR21 U2300 ( .A(n2845), .B(n2893), .Q(n3052) );
  OAI221 U2301 ( .A(n3053), .B(n2891), .C(n3054), .D(n2985), .Q(n1939) );
  XNR21 U2302 ( .A(n2846), .B(n2893), .Q(n3053) );
  OAI221 U2303 ( .A(n3054), .B(n2891), .C(n3055), .D(n2985), .Q(n1938) );
  XNR21 U2304 ( .A(n2847), .B(n2893), .Q(n3054) );
  AOI211 U2305 ( .A(n2985), .B(n2756), .C(n3055), .Q(n3056) );
  XNR21 U2306 ( .A(n2848), .B(n2893), .Q(n3055) );
  NOR22 U2307 ( .A(n2817), .B(n2986), .Q(n1936) );
  XNR21 U2308 ( .A(n2986), .B(n2897), .Q(n3057) );
  OAI221 U2309 ( .A(n3058), .B(n2997), .C(n2817), .D(n3059), .Q(n1934) );
  XNR21 U2310 ( .A(n2818), .B(n2895), .Q(n3058) );
  OAI221 U2311 ( .A(n3059), .B(n2858), .C(n2816), .D(n3060), .Q(n1933) );
  XNR21 U2312 ( .A(n2819), .B(n2895), .Q(n3059) );
  XNR21 U2313 ( .A(n2820), .B(n2895), .Q(n3060) );
  OAI221 U2314 ( .A(n3061), .B(n2857), .C(n2816), .D(n3062), .Q(n1931) );
  XNR21 U2315 ( .A(n2821), .B(n2895), .Q(n3061) );
  OAI221 U2316 ( .A(n3062), .B(n2858), .C(n2816), .D(n3063), .Q(n1930) );
  XNR21 U2317 ( .A(n2822), .B(n2895), .Q(n3062) );
  OAI221 U2318 ( .A(n3063), .B(n2857), .C(n2816), .D(n3064), .Q(n1929) );
  XNR21 U2319 ( .A(n2823), .B(n2895), .Q(n3063) );
  OAI221 U2320 ( .A(n3064), .B(n2857), .C(n2816), .D(n3065), .Q(n1928) );
  XNR21 U2321 ( .A(n2824), .B(n2895), .Q(n3064) );
  OAI221 U2322 ( .A(n3065), .B(n2857), .C(n2816), .D(n3066), .Q(n1927) );
  XNR21 U2323 ( .A(n2825), .B(n2895), .Q(n3065) );
  OAI221 U2324 ( .A(n3066), .B(n2857), .C(n2816), .D(n3067), .Q(n1926) );
  XNR21 U2325 ( .A(n2826), .B(n2895), .Q(n3066) );
  OAI221 U2326 ( .A(n3067), .B(n2857), .C(n2816), .D(n3068), .Q(n1925) );
  XNR21 U2327 ( .A(n2827), .B(n2896), .Q(n3067) );
  OAI221 U2328 ( .A(n3068), .B(n2857), .C(n2816), .D(n3069), .Q(n1924) );
  XNR21 U2329 ( .A(n2828), .B(n2896), .Q(n3068) );
  OAI221 U2330 ( .A(n3069), .B(n2857), .C(n2816), .D(n3070), .Q(n1923) );
  XNR21 U2331 ( .A(n2829), .B(n2896), .Q(n3069) );
  OAI221 U2332 ( .A(n3070), .B(n2858), .C(n2816), .D(n3071), .Q(n1922) );
  XNR21 U2333 ( .A(n2830), .B(n2896), .Q(n3070) );
  OAI221 U2334 ( .A(n3071), .B(n2858), .C(n2816), .D(n3072), .Q(n1921) );
  XNR21 U2335 ( .A(n2831), .B(n2896), .Q(n3071) );
  OAI221 U2336 ( .A(n3072), .B(n2858), .C(n2816), .D(n3073), .Q(n1920) );
  XNR21 U2337 ( .A(n2832), .B(n2896), .Q(n3072) );
  OAI221 U2338 ( .A(n3073), .B(n2858), .C(n2816), .D(n3074), .Q(n1919) );
  XNR21 U2339 ( .A(n2833), .B(n2896), .Q(n3073) );
  OAI221 U2340 ( .A(n3074), .B(n2858), .C(n2816), .D(n3075), .Q(n1918) );
  XNR21 U2341 ( .A(n2834), .B(n2896), .Q(n3074) );
  OAI221 U2342 ( .A(n3075), .B(n2858), .C(n2816), .D(n3076), .Q(n1917) );
  XNR21 U2343 ( .A(n2835), .B(n2896), .Q(n3075) );
  OAI221 U2344 ( .A(n3076), .B(n2858), .C(n2816), .D(n3077), .Q(n1916) );
  XNR21 U2345 ( .A(n2836), .B(n2896), .Q(n3076) );
  OAI221 U2346 ( .A(n3077), .B(n2858), .C(n2816), .D(n3078), .Q(n1915) );
  XNR21 U2347 ( .A(n2837), .B(n2896), .Q(n3077) );
  OAI221 U2348 ( .A(n3078), .B(n2858), .C(n2816), .D(n3079), .Q(n1914) );
  XNR21 U2349 ( .A(n2838), .B(n2896), .Q(n3078) );
  OAI221 U2350 ( .A(n3079), .B(n2858), .C(n2816), .D(n3080), .Q(n1913) );
  XNR21 U2351 ( .A(n2839), .B(n2896), .Q(n3079) );
  OAI221 U2352 ( .A(n3080), .B(n2858), .C(n2816), .D(n3081), .Q(n1912) );
  XNR21 U2353 ( .A(n2840), .B(n2896), .Q(n3080) );
  OAI221 U2354 ( .A(n3081), .B(n2858), .C(n2816), .D(n3082), .Q(n1911) );
  XNR21 U2355 ( .A(n2841), .B(n2896), .Q(n3081) );
  OAI221 U2356 ( .A(n3082), .B(n2857), .C(n2816), .D(n3083), .Q(n1910) );
  XNR21 U2357 ( .A(n2842), .B(n2896), .Q(n3082) );
  OAI221 U2358 ( .A(n3083), .B(n2858), .C(n2816), .D(n3084), .Q(n1909) );
  XNR21 U2359 ( .A(n2843), .B(n2896), .Q(n3083) );
  OAI221 U2360 ( .A(n3084), .B(n2857), .C(n2816), .D(n3085), .Q(n1908) );
  XNR21 U2361 ( .A(n2844), .B(n2896), .Q(n3084) );
  OAI221 U2362 ( .A(n3085), .B(n2857), .C(n2816), .D(n3086), .Q(n1907) );
  XNR21 U2363 ( .A(n2845), .B(n2896), .Q(n3085) );
  OAI221 U2364 ( .A(n3086), .B(n2858), .C(n2816), .D(n2996), .Q(n1906) );
  XNR21 U2365 ( .A(n2847), .B(n2896), .Q(n2996) );
  XNR21 U2366 ( .A(n2846), .B(n2896), .Q(n3086) );
  AOI211 U2367 ( .A(n2857), .B(n2816), .C(n2757), .Q(n3087) );
  NOR22 U2368 ( .A(n2814), .B(n2850), .Q(n1904) );
  XNR21 U2369 ( .A(n2818), .B(n2898), .Q(n3089) );
  OAI221 U2370 ( .A(n3090), .B(n2999), .C(n2814), .D(n3091), .Q(n1901) );
  XNR21 U2371 ( .A(n2819), .B(n2898), .Q(n3090) );
  XNR21 U2372 ( .A(n2820), .B(n2898), .Q(n3091) );
  OAI221 U2373 ( .A(n3092), .B(n2859), .C(n2814), .D(n3093), .Q(n1899) );
  XNR21 U2374 ( .A(n2821), .B(n2898), .Q(n3092) );
  OAI221 U2375 ( .A(n3093), .B(n2860), .C(n2814), .D(n3094), .Q(n1898) );
  XNR21 U2376 ( .A(n2822), .B(n2898), .Q(n3093) );
  OAI221 U2377 ( .A(n3094), .B(n2860), .C(n2814), .D(n3095), .Q(n1897) );
  XNR21 U2378 ( .A(n2823), .B(n2898), .Q(n3094) );
  OAI221 U2379 ( .A(n3095), .B(n2860), .C(n2814), .D(n3096), .Q(n1896) );
  XNR21 U2380 ( .A(n2824), .B(n2898), .Q(n3095) );
  OAI221 U2381 ( .A(n3096), .B(n2860), .C(n2814), .D(n3097), .Q(n1895) );
  XNR21 U2382 ( .A(n2825), .B(n2898), .Q(n3096) );
  OAI221 U2383 ( .A(n3097), .B(n2860), .C(n2814), .D(n3098), .Q(n1894) );
  XNR21 U2384 ( .A(n2826), .B(n2898), .Q(n3097) );
  OAI221 U2385 ( .A(n3098), .B(n2860), .C(n2814), .D(n3099), .Q(n1893) );
  XNR21 U2386 ( .A(n2827), .B(n2899), .Q(n3098) );
  OAI221 U2387 ( .A(n3099), .B(n2860), .C(n2814), .D(n3100), .Q(n1892) );
  XNR21 U2388 ( .A(n2828), .B(n2899), .Q(n3099) );
  OAI221 U2389 ( .A(n3100), .B(n2860), .C(n2814), .D(n3101), .Q(n1891) );
  XNR21 U2390 ( .A(n2829), .B(n2899), .Q(n3100) );
  OAI221 U2391 ( .A(n3101), .B(n2859), .C(n2814), .D(n3102), .Q(n1890) );
  XNR21 U2392 ( .A(n2830), .B(n2899), .Q(n3101) );
  OAI221 U2393 ( .A(n3102), .B(n2859), .C(n2814), .D(n3103), .Q(n1889) );
  XNR21 U2394 ( .A(n2831), .B(n2899), .Q(n3102) );
  OAI221 U2395 ( .A(n3103), .B(n2859), .C(n2815), .D(n3104), .Q(n1888) );
  XNR21 U2396 ( .A(n2832), .B(n2899), .Q(n3103) );
  OAI221 U2397 ( .A(n3104), .B(n2859), .C(n2815), .D(n3105), .Q(n1887) );
  XNR21 U2398 ( .A(n2833), .B(n2899), .Q(n3104) );
  OAI221 U2399 ( .A(n3105), .B(n2859), .C(n2815), .D(n3106), .Q(n1886) );
  XNR21 U2400 ( .A(n2834), .B(n2899), .Q(n3105) );
  OAI221 U2401 ( .A(n3106), .B(n2859), .C(n2815), .D(n3107), .Q(n1885) );
  XNR21 U2402 ( .A(n2835), .B(n2899), .Q(n3106) );
  OAI221 U2403 ( .A(n3107), .B(n2860), .C(n2815), .D(n3108), .Q(n1884) );
  XNR21 U2404 ( .A(n2836), .B(n2899), .Q(n3107) );
  OAI221 U2405 ( .A(n3108), .B(n2860), .C(n2815), .D(n3109), .Q(n1883) );
  XNR21 U2406 ( .A(n2837), .B(n2899), .Q(n3108) );
  OAI221 U2407 ( .A(n3109), .B(n2860), .C(n2815), .D(n3110), .Q(n1882) );
  XNR21 U2408 ( .A(n2838), .B(n2899), .Q(n3109) );
  OAI221 U2409 ( .A(n3110), .B(n2860), .C(n2815), .D(n3111), .Q(n1881) );
  XNR21 U2410 ( .A(n2839), .B(n2899), .Q(n3110) );
  OAI221 U2411 ( .A(n3111), .B(n2860), .C(n2815), .D(n3112), .Q(n1880) );
  XNR21 U2412 ( .A(n2840), .B(n2899), .Q(n3111) );
  OAI221 U2413 ( .A(n3112), .B(n2860), .C(n2815), .D(n3113), .Q(n1879) );
  XNR21 U2414 ( .A(n2841), .B(n2899), .Q(n3112) );
  OAI221 U2415 ( .A(n3113), .B(n2860), .C(n2815), .D(n3114), .Q(n1878) );
  XNR21 U2416 ( .A(n2842), .B(n2899), .Q(n3113) );
  OAI221 U2417 ( .A(n3114), .B(n2860), .C(n2815), .D(n3115), .Q(n1877) );
  XNR21 U2418 ( .A(n2843), .B(n2899), .Q(n3114) );
  OAI221 U2419 ( .A(n3115), .B(n2860), .C(n2815), .D(n3116), .Q(n1876) );
  XNR21 U2420 ( .A(n2844), .B(n2899), .Q(n3115) );
  OAI221 U2421 ( .A(n3116), .B(n2860), .C(n2815), .D(n3117), .Q(n1875) );
  XNR21 U2422 ( .A(n2845), .B(n2899), .Q(n3116) );
  OAI221 U2423 ( .A(n3117), .B(n2860), .C(n2815), .D(n2998), .Q(n1874) );
  XNR21 U2424 ( .A(n2847), .B(n2899), .Q(n2998) );
  XNR21 U2425 ( .A(n2846), .B(n2899), .Q(n3117) );
  AOI211 U2426 ( .A(n2860), .B(n2815), .C(n2753), .Q(n3118) );
  OAI221 U2427 ( .A(n3119), .B(n3001), .C(n2813), .D(n3120), .Q(n1871) );
  XNR21 U2428 ( .A(n2850), .B(n2903), .Q(n3119) );
  OAI221 U2429 ( .A(n3120), .B(n3001), .C(n2813), .D(n3121), .Q(n1870) );
  XNR21 U2430 ( .A(n2818), .B(n2901), .Q(n3120) );
  OAI221 U2431 ( .A(n3121), .B(n3001), .C(n2813), .D(n3122), .Q(n1869) );
  XNR21 U2432 ( .A(n2819), .B(n2901), .Q(n3121) );
  OAI221 U2433 ( .A(n3122), .B(n2861), .C(n2813), .D(n3123), .Q(n1868) );
  XNR21 U2434 ( .A(n2820), .B(n2901), .Q(n3122) );
  OAI221 U2435 ( .A(n3123), .B(n2861), .C(n2813), .D(n3124), .Q(n1867) );
  XNR21 U2436 ( .A(n2821), .B(n2901), .Q(n3123) );
  OAI221 U2437 ( .A(n3124), .B(n2861), .C(n2813), .D(n3125), .Q(n1866) );
  XNR21 U2438 ( .A(n2822), .B(n2901), .Q(n3124) );
  OAI221 U2439 ( .A(n3125), .B(n2861), .C(n2813), .D(n3126), .Q(n1865) );
  XNR21 U2440 ( .A(n2823), .B(n2901), .Q(n3125) );
  OAI221 U2441 ( .A(n3126), .B(n2861), .C(n2813), .D(n3127), .Q(n1864) );
  XNR21 U2442 ( .A(n2824), .B(n2901), .Q(n3126) );
  OAI221 U2443 ( .A(n3127), .B(n2861), .C(n2813), .D(n3128), .Q(n1863) );
  XNR21 U2444 ( .A(n2825), .B(n2901), .Q(n3127) );
  OAI221 U2445 ( .A(n3128), .B(n2861), .C(n2813), .D(n3129), .Q(n1862) );
  XNR21 U2446 ( .A(n2826), .B(n2901), .Q(n3128) );
  OAI221 U2447 ( .A(n3129), .B(n2861), .C(n2813), .D(n3130), .Q(n1861) );
  XNR21 U2448 ( .A(n2827), .B(n2902), .Q(n3129) );
  OAI221 U2449 ( .A(n3130), .B(n2861), .C(n2813), .D(n3131), .Q(n1860) );
  XNR21 U2450 ( .A(n2828), .B(n2902), .Q(n3130) );
  OAI221 U2451 ( .A(n3131), .B(n2861), .C(n2813), .D(n3132), .Q(n1859) );
  XNR21 U2452 ( .A(n2829), .B(n2902), .Q(n3131) );
  OAI221 U2453 ( .A(n3132), .B(n2861), .C(n2813), .D(n3133), .Q(n1858) );
  XNR21 U2454 ( .A(n2830), .B(n2902), .Q(n3132) );
  OAI221 U2455 ( .A(n3133), .B(n2861), .C(n2813), .D(n3134), .Q(n1857) );
  XNR21 U2456 ( .A(n2831), .B(n2902), .Q(n3133) );
  OAI221 U2457 ( .A(n3134), .B(n2861), .C(n2977), .D(n3135), .Q(n1856) );
  XNR21 U2458 ( .A(n2832), .B(n2902), .Q(n3134) );
  OAI221 U2459 ( .A(n3135), .B(n2861), .C(n2977), .D(n3136), .Q(n1855) );
  XNR21 U2460 ( .A(n2833), .B(n2902), .Q(n3135) );
  OAI221 U2461 ( .A(n3136), .B(n2861), .C(n2977), .D(n3137), .Q(n1854) );
  XNR21 U2462 ( .A(n2834), .B(n2902), .Q(n3136) );
  OAI221 U2463 ( .A(n3137), .B(n2861), .C(n2977), .D(n3138), .Q(n1853) );
  XNR21 U2464 ( .A(n2835), .B(n2902), .Q(n3137) );
  OAI221 U2465 ( .A(n3138), .B(n2861), .C(n2977), .D(n3139), .Q(n1852) );
  XNR21 U2466 ( .A(n2836), .B(n2902), .Q(n3138) );
  OAI221 U2467 ( .A(n3139), .B(n2861), .C(n2977), .D(n3140), .Q(n1851) );
  XNR21 U2468 ( .A(n2837), .B(n2902), .Q(n3139) );
  OAI221 U2469 ( .A(n3140), .B(n2861), .C(n2977), .D(n3141), .Q(n1850) );
  XNR21 U2470 ( .A(n2838), .B(n2902), .Q(n3140) );
  OAI221 U2471 ( .A(n3141), .B(n2861), .C(n2977), .D(n3142), .Q(n1849) );
  XNR21 U2472 ( .A(n2839), .B(n2902), .Q(n3141) );
  OAI221 U2473 ( .A(n3142), .B(n2861), .C(n2977), .D(n3143), .Q(n1848) );
  XNR21 U2474 ( .A(n2840), .B(n2902), .Q(n3142) );
  OAI221 U2475 ( .A(n3143), .B(n2861), .C(n2977), .D(n3144), .Q(n1847) );
  XNR21 U2476 ( .A(n2841), .B(n2902), .Q(n3143) );
  OAI221 U2477 ( .A(n3144), .B(n2861), .C(n2977), .D(n3145), .Q(n1846) );
  XNR21 U2478 ( .A(n2842), .B(n2902), .Q(n3144) );
  OAI221 U2479 ( .A(n3145), .B(n2861), .C(n2977), .D(n3146), .Q(n1845) );
  XNR21 U2480 ( .A(n2843), .B(n2902), .Q(n3145) );
  OAI221 U2481 ( .A(n3146), .B(n2861), .C(n2977), .D(n3147), .Q(n1844) );
  XNR21 U2482 ( .A(n2844), .B(n2902), .Q(n3146) );
  OAI221 U2483 ( .A(n3147), .B(n2861), .C(n2977), .D(n3148), .Q(n1843) );
  XNR21 U2484 ( .A(n2845), .B(n2902), .Q(n3147) );
  OAI221 U2485 ( .A(n3148), .B(n2861), .C(n2977), .D(n3000), .Q(n1842) );
  XNR21 U2486 ( .A(n2847), .B(n2902), .Q(n3000) );
  XNR21 U2487 ( .A(n2846), .B(n2902), .Q(n3148) );
  AOI211 U2488 ( .A(n2861), .B(n2977), .C(n2754), .Q(n3149) );
  NOR22 U2489 ( .A(n2974), .B(n2849), .Q(n1840) );
  OAI221 U2490 ( .A(n3150), .B(n3003), .C(n2974), .D(n3151), .Q(n1839) );
  XNR21 U2491 ( .A(n2849), .B(n2906), .Q(n3150) );
  OAI221 U2492 ( .A(n3151), .B(n3003), .C(n2974), .D(n3152), .Q(n1838) );
  XNR21 U2493 ( .A(n2818), .B(n2904), .Q(n3151) );
  OAI221 U2494 ( .A(n3152), .B(n2862), .C(n2974), .D(n3153), .Q(n1837) );
  XNR21 U2495 ( .A(n2819), .B(n2904), .Q(n3152) );
  OAI221 U2496 ( .A(n3153), .B(n2862), .C(n2974), .D(n3154), .Q(n1836) );
  XNR21 U2497 ( .A(n2820), .B(n2904), .Q(n3153) );
  OAI221 U2498 ( .A(n3154), .B(n2862), .C(n2974), .D(n3155), .Q(n1835) );
  XNR21 U2499 ( .A(n2821), .B(n2904), .Q(n3154) );
  OAI221 U2500 ( .A(n3155), .B(n2862), .C(n2974), .D(n3156), .Q(n1834) );
  XNR21 U2501 ( .A(n2822), .B(n2904), .Q(n3155) );
  OAI221 U2502 ( .A(n3156), .B(n2862), .C(n2974), .D(n3157), .Q(n1833) );
  XNR21 U2503 ( .A(n2823), .B(n2904), .Q(n3156) );
  OAI221 U2504 ( .A(n3157), .B(n2862), .C(n2974), .D(n3158), .Q(n1832) );
  XNR21 U2505 ( .A(n2824), .B(n2904), .Q(n3157) );
  OAI221 U2506 ( .A(n3158), .B(n2862), .C(n2974), .D(n3159), .Q(n1831) );
  XNR21 U2507 ( .A(n2825), .B(n2904), .Q(n3158) );
  OAI221 U2508 ( .A(n3159), .B(n2862), .C(n2974), .D(n3160), .Q(n1830) );
  XNR21 U2509 ( .A(n2826), .B(n2904), .Q(n3159) );
  OAI221 U2510 ( .A(n3160), .B(n2862), .C(n2974), .D(n3161), .Q(n1829) );
  XNR21 U2511 ( .A(n2827), .B(n2905), .Q(n3160) );
  OAI221 U2512 ( .A(n3161), .B(n2862), .C(n2974), .D(n3162), .Q(n1828) );
  XNR21 U2513 ( .A(n2828), .B(n2905), .Q(n3161) );
  OAI221 U2514 ( .A(n3162), .B(n2862), .C(n2974), .D(n3163), .Q(n1827) );
  XNR21 U2515 ( .A(n2829), .B(n2905), .Q(n3162) );
  OAI221 U2516 ( .A(n3163), .B(n2862), .C(n2974), .D(n3164), .Q(n1826) );
  XNR21 U2517 ( .A(n2830), .B(n2905), .Q(n3163) );
  OAI221 U2518 ( .A(n3164), .B(n2862), .C(n2974), .D(n3165), .Q(n1825) );
  XNR21 U2519 ( .A(n2831), .B(n2905), .Q(n3164) );
  OAI221 U2520 ( .A(n3165), .B(n2862), .C(n2974), .D(n3166), .Q(n1824) );
  XNR21 U2521 ( .A(n2832), .B(n2905), .Q(n3165) );
  OAI221 U2522 ( .A(n3166), .B(n2862), .C(n2974), .D(n3167), .Q(n1823) );
  XNR21 U2523 ( .A(n2833), .B(n2905), .Q(n3166) );
  OAI221 U2524 ( .A(n3167), .B(n2862), .C(n2974), .D(n3168), .Q(n1822) );
  XNR21 U2525 ( .A(n2834), .B(n2905), .Q(n3167) );
  OAI221 U2526 ( .A(n3168), .B(n2862), .C(n2974), .D(n3169), .Q(n1821) );
  XNR21 U2527 ( .A(n2835), .B(n2905), .Q(n3168) );
  OAI221 U2528 ( .A(n3169), .B(n2862), .C(n2974), .D(n3170), .Q(n1820) );
  XNR21 U2529 ( .A(n2836), .B(n2905), .Q(n3169) );
  OAI221 U2530 ( .A(n3170), .B(n2862), .C(n2974), .D(n3171), .Q(n1819) );
  XNR21 U2531 ( .A(n2837), .B(n2905), .Q(n3170) );
  OAI221 U2532 ( .A(n3171), .B(n2862), .C(n2974), .D(n3172), .Q(n1818) );
  XNR21 U2533 ( .A(n2838), .B(n2905), .Q(n3171) );
  OAI221 U2534 ( .A(n3172), .B(n2862), .C(n2974), .D(n3173), .Q(n1817) );
  XNR21 U2535 ( .A(n2839), .B(n2905), .Q(n3172) );
  OAI221 U2536 ( .A(n3173), .B(n2862), .C(n2974), .D(n3174), .Q(n1816) );
  XNR21 U2537 ( .A(n2840), .B(n2905), .Q(n3173) );
  OAI221 U2538 ( .A(n3174), .B(n2862), .C(n2974), .D(n3175), .Q(n1815) );
  XNR21 U2539 ( .A(n2841), .B(n2905), .Q(n3174) );
  OAI221 U2540 ( .A(n3175), .B(n2862), .C(n2974), .D(n3176), .Q(n1814) );
  XNR21 U2541 ( .A(n2842), .B(n2905), .Q(n3175) );
  OAI221 U2542 ( .A(n3176), .B(n2862), .C(n2974), .D(n3177), .Q(n1813) );
  XNR21 U2543 ( .A(n2843), .B(n2905), .Q(n3176) );
  OAI221 U2544 ( .A(n3177), .B(n2862), .C(n2974), .D(n3178), .Q(n1812) );
  XNR21 U2545 ( .A(n2844), .B(n2905), .Q(n3177) );
  OAI221 U2546 ( .A(n3178), .B(n2862), .C(n2974), .D(n3179), .Q(n1811) );
  XNR21 U2547 ( .A(n2845), .B(n2905), .Q(n3178) );
  OAI221 U2548 ( .A(n3179), .B(n2862), .C(n2974), .D(n3002), .Q(n1810) );
  XNR21 U2549 ( .A(n2847), .B(n2905), .Q(n3002) );
  XNR21 U2550 ( .A(n2846), .B(n2905), .Q(n3179) );
  AOI211 U2551 ( .A(n2862), .B(n2974), .C(n2755), .Q(n3180) );
  NOR22 U2552 ( .A(n2971), .B(n2986), .Q(n1808) );
  OAI221 U2553 ( .A(n3181), .B(n3005), .C(n2971), .D(n3182), .Q(n1807) );
  XNR21 U2554 ( .A(n2849), .B(n2908), .Q(n3181) );
  OAI221 U2555 ( .A(n3182), .B(n3005), .C(n2971), .D(n3183), .Q(n1806) );
  XNR21 U2556 ( .A(n2818), .B(n2907), .Q(n3182) );
  OAI221 U2557 ( .A(n3183), .B(n2863), .C(n2971), .D(n3184), .Q(n1805) );
  XNR21 U2558 ( .A(n2819), .B(n2907), .Q(n3183) );
  OAI221 U2559 ( .A(n3184), .B(n2863), .C(n2971), .D(n3185), .Q(n1804) );
  XNR21 U2560 ( .A(n2820), .B(n2907), .Q(n3184) );
  OAI221 U2561 ( .A(n3185), .B(n2863), .C(n2971), .D(n3186), .Q(n1803) );
  XNR21 U2562 ( .A(n2821), .B(n2907), .Q(n3185) );
  OAI221 U2563 ( .A(n3186), .B(n2863), .C(n2971), .D(n3187), .Q(n1802) );
  XNR21 U2564 ( .A(n2822), .B(n2907), .Q(n3186) );
  OAI221 U2565 ( .A(n3187), .B(n2863), .C(n2971), .D(n3188), .Q(n1801) );
  XNR21 U2566 ( .A(n2823), .B(n2907), .Q(n3187) );
  OAI221 U2567 ( .A(n3188), .B(n2863), .C(n2971), .D(n3189), .Q(n1800) );
  XNR21 U2568 ( .A(n2824), .B(n2907), .Q(n3188) );
  OAI221 U2569 ( .A(n3189), .B(n2863), .C(n2971), .D(n3190), .Q(n1799) );
  XNR21 U2570 ( .A(n2825), .B(n2907), .Q(n3189) );
  OAI221 U2571 ( .A(n3190), .B(n2863), .C(n2971), .D(n3191), .Q(n1798) );
  XNR21 U2572 ( .A(n2826), .B(n2907), .Q(n3190) );
  OAI221 U2573 ( .A(n3191), .B(n2863), .C(n2971), .D(n3192), .Q(n1797) );
  XNR21 U2574 ( .A(n2827), .B(n2907), .Q(n3191) );
  OAI221 U2575 ( .A(n3192), .B(n2863), .C(n2971), .D(n3193), .Q(n1796) );
  XNR21 U2576 ( .A(n2828), .B(n2907), .Q(n3192) );
  OAI221 U2577 ( .A(n3193), .B(n2863), .C(n2971), .D(n3194), .Q(n1795) );
  XNR21 U2578 ( .A(n2829), .B(n2907), .Q(n3193) );
  OAI221 U2579 ( .A(n3194), .B(n2863), .C(n2971), .D(n3195), .Q(n1794) );
  XNR21 U2580 ( .A(n2830), .B(n2907), .Q(n3194) );
  OAI221 U2581 ( .A(n3195), .B(n2863), .C(n2971), .D(n3196), .Q(n1793) );
  XNR21 U2582 ( .A(n2831), .B(n2907), .Q(n3195) );
  OAI221 U2583 ( .A(n3196), .B(n2863), .C(n2971), .D(n3197), .Q(n1792) );
  XNR21 U2584 ( .A(n2832), .B(n2907), .Q(n3196) );
  OAI221 U2585 ( .A(n3197), .B(n2863), .C(n2971), .D(n3198), .Q(n1791) );
  XNR21 U2586 ( .A(n2833), .B(n2907), .Q(n3197) );
  OAI221 U2587 ( .A(n3198), .B(n2863), .C(n2971), .D(n3199), .Q(n1790) );
  XNR21 U2588 ( .A(n2834), .B(n2907), .Q(n3198) );
  OAI221 U2589 ( .A(n3199), .B(n2863), .C(n2971), .D(n3200), .Q(n1789) );
  XNR21 U2590 ( .A(n2835), .B(n2907), .Q(n3199) );
  OAI221 U2591 ( .A(n3200), .B(n2863), .C(n2971), .D(n3201), .Q(n1788) );
  XNR21 U2592 ( .A(n2836), .B(n2907), .Q(n3200) );
  OAI221 U2593 ( .A(n3201), .B(n2863), .C(n2971), .D(n3202), .Q(n1787) );
  XNR21 U2594 ( .A(n2837), .B(n2907), .Q(n3201) );
  OAI221 U2595 ( .A(n3202), .B(n2863), .C(n2971), .D(n3203), .Q(n1786) );
  XNR21 U2596 ( .A(n2838), .B(n2907), .Q(n3202) );
  OAI221 U2597 ( .A(n3203), .B(n2863), .C(n2971), .D(n3204), .Q(n1785) );
  XNR21 U2598 ( .A(n2839), .B(n2907), .Q(n3203) );
  OAI221 U2599 ( .A(n3204), .B(n2863), .C(n2971), .D(n3205), .Q(n1784) );
  XNR21 U2600 ( .A(n2840), .B(n2907), .Q(n3204) );
  OAI221 U2601 ( .A(n3205), .B(n2863), .C(n2971), .D(n3206), .Q(n1783) );
  XNR21 U2602 ( .A(n2841), .B(n2907), .Q(n3205) );
  OAI221 U2603 ( .A(n3206), .B(n2863), .C(n2971), .D(n3207), .Q(n1782) );
  XNR21 U2604 ( .A(n2842), .B(a[11]), .Q(n3206) );
  OAI221 U2605 ( .A(n3207), .B(n2863), .C(n2971), .D(n3208), .Q(n1781) );
  XNR21 U2606 ( .A(n2843), .B(a[11]), .Q(n3207) );
  OAI221 U2607 ( .A(n3208), .B(n2863), .C(n2971), .D(n3209), .Q(n1780) );
  XNR21 U2608 ( .A(n2844), .B(a[11]), .Q(n3208) );
  OAI221 U2609 ( .A(n3209), .B(n2863), .C(n2971), .D(n3210), .Q(n1779) );
  XNR21 U2610 ( .A(n2845), .B(a[11]), .Q(n3209) );
  OAI221 U2611 ( .A(n3210), .B(n2863), .C(n2971), .D(n3004), .Q(n1778) );
  XNR21 U2612 ( .A(n2847), .B(a[11]), .Q(n3004) );
  XNR21 U2613 ( .A(n2846), .B(a[11]), .Q(n3210) );
  AOI211 U2614 ( .A(n2863), .B(n2971), .C(n2739), .Q(n3211) );
  NOR22 U2615 ( .A(n2968), .B(n2986), .Q(n1776) );
  OAI221 U2616 ( .A(n3212), .B(n2994), .C(n2968), .D(n3213), .Q(n1775) );
  XNR21 U2617 ( .A(n2849), .B(n2910), .Q(n3212) );
  XNR21 U2618 ( .A(n2818), .B(n2909), .Q(n3213) );
  OAI221 U2619 ( .A(n3214), .B(n2856), .C(n2968), .D(n3215), .Q(n1773) );
  XNR21 U2620 ( .A(n2819), .B(n2909), .Q(n3214) );
  OAI221 U2621 ( .A(n3215), .B(n2856), .C(n2968), .D(n3216), .Q(n1772) );
  XNR21 U2622 ( .A(n2820), .B(n2909), .Q(n3215) );
  OAI221 U2623 ( .A(n3216), .B(n2856), .C(n2968), .D(n3217), .Q(n1771) );
  XNR21 U2624 ( .A(n2821), .B(n2909), .Q(n3216) );
  OAI221 U2625 ( .A(n3217), .B(n2856), .C(n2968), .D(n3218), .Q(n1770) );
  XNR21 U2626 ( .A(n2822), .B(n2909), .Q(n3217) );
  OAI221 U2627 ( .A(n3218), .B(n2856), .C(n2968), .D(n3219), .Q(n1769) );
  XNR21 U2628 ( .A(n2823), .B(n2909), .Q(n3218) );
  OAI221 U2629 ( .A(n3219), .B(n2856), .C(n2968), .D(n3220), .Q(n1768) );
  XNR21 U2630 ( .A(n2824), .B(n2909), .Q(n3219) );
  OAI221 U2631 ( .A(n3220), .B(n2856), .C(n2968), .D(n3221), .Q(n1767) );
  XNR21 U2632 ( .A(n2825), .B(n2909), .Q(n3220) );
  OAI221 U2633 ( .A(n3221), .B(n2856), .C(n2968), .D(n3222), .Q(n1766) );
  XNR21 U2634 ( .A(n2826), .B(n2909), .Q(n3221) );
  OAI221 U2635 ( .A(n3222), .B(n2856), .C(n2968), .D(n3223), .Q(n1765) );
  XNR21 U2636 ( .A(n2827), .B(n2909), .Q(n3222) );
  OAI221 U2637 ( .A(n3223), .B(n2856), .C(n2968), .D(n3224), .Q(n1764) );
  XNR21 U2638 ( .A(n2828), .B(n2909), .Q(n3223) );
  OAI221 U2639 ( .A(n3224), .B(n2856), .C(n2968), .D(n3225), .Q(n1763) );
  XNR21 U2640 ( .A(n2829), .B(n2909), .Q(n3224) );
  OAI221 U2641 ( .A(n3225), .B(n2856), .C(n2968), .D(n3226), .Q(n1762) );
  XNR21 U2642 ( .A(n2830), .B(n2909), .Q(n3225) );
  OAI221 U2643 ( .A(n3226), .B(n2856), .C(n2968), .D(n3227), .Q(n1761) );
  XNR21 U2644 ( .A(n2831), .B(n2909), .Q(n3226) );
  OAI221 U2645 ( .A(n3227), .B(n2856), .C(n2968), .D(n3228), .Q(n1760) );
  XNR21 U2646 ( .A(n2832), .B(n2909), .Q(n3227) );
  OAI221 U2647 ( .A(n3228), .B(n2856), .C(n2968), .D(n3229), .Q(n1759) );
  XNR21 U2648 ( .A(n2833), .B(n2909), .Q(n3228) );
  OAI221 U2649 ( .A(n3229), .B(n2856), .C(n2968), .D(n3230), .Q(n1758) );
  XNR21 U2650 ( .A(n2834), .B(n2909), .Q(n3229) );
  OAI221 U2651 ( .A(n3230), .B(n2856), .C(n2968), .D(n2993), .Q(n1757) );
  XNR21 U2652 ( .A(n2836), .B(n2909), .Q(n2993) );
  XNR21 U2653 ( .A(n2835), .B(n2909), .Q(n3230) );
  OAI221 U2654 ( .A(n2995), .B(n2856), .C(n2968), .D(n3231), .Q(n1755) );
  XNR21 U2655 ( .A(n2837), .B(n2909), .Q(n2995) );
  OAI221 U2656 ( .A(n3231), .B(n2856), .C(n2968), .D(n3232), .Q(n1754) );
  XNR21 U2657 ( .A(n2838), .B(n2909), .Q(n3231) );
  OAI221 U2658 ( .A(n3232), .B(n2856), .C(n2968), .D(n3233), .Q(n1753) );
  XNR21 U2659 ( .A(n2839), .B(n2909), .Q(n3232) );
  OAI221 U2660 ( .A(n3233), .B(n2856), .C(n2968), .D(n3234), .Q(n1752) );
  XNR21 U2661 ( .A(n2840), .B(n2909), .Q(n3233) );
  OAI221 U2662 ( .A(n3234), .B(n2856), .C(n2968), .D(n3235), .Q(n1751) );
  XNR21 U2663 ( .A(n2841), .B(n2909), .Q(n3234) );
  OAI221 U2664 ( .A(n3235), .B(n2856), .C(n2968), .D(n3236), .Q(n1750) );
  XNR21 U2665 ( .A(n2842), .B(n2909), .Q(n3235) );
  OAI221 U2666 ( .A(n3236), .B(n2856), .C(n2968), .D(n3237), .Q(n1749) );
  XNR21 U2667 ( .A(n2843), .B(n2909), .Q(n3236) );
  OAI221 U2668 ( .A(n3237), .B(n2856), .C(n2968), .D(n3238), .Q(n1748) );
  XNR21 U2669 ( .A(n2844), .B(n2909), .Q(n3237) );
  OAI221 U2670 ( .A(n3238), .B(n2856), .C(n2968), .D(n3239), .Q(n1747) );
  XNR21 U2671 ( .A(n2845), .B(a[13]), .Q(n3238) );
  OAI221 U2672 ( .A(n3239), .B(n2856), .C(n2968), .D(n3006), .Q(n1746) );
  XNR21 U2673 ( .A(n2847), .B(a[13]), .Q(n3006) );
  XNR21 U2674 ( .A(n2846), .B(a[13]), .Q(n3239) );
  AOI211 U2675 ( .A(n2856), .B(n2968), .C(n2740), .Q(n3240) );
  NOR22 U2676 ( .A(n2965), .B(n2986), .Q(n1744) );
  OAI221 U2677 ( .A(n3241), .B(n3008), .C(n2965), .D(n3242), .Q(n1743) );
  XNR21 U2678 ( .A(n2849), .B(n2913), .Q(n3241) );
  OAI221 U2679 ( .A(n3242), .B(n2864), .C(n2965), .D(n3243), .Q(n1742) );
  XNR21 U2680 ( .A(n2818), .B(n2911), .Q(n3242) );
  OAI221 U2681 ( .A(n3243), .B(n2864), .C(n2965), .D(n3244), .Q(n1741) );
  XNR21 U2682 ( .A(n2819), .B(n2911), .Q(n3243) );
  OAI221 U2683 ( .A(n3244), .B(n2864), .C(n2965), .D(n3245), .Q(n1740) );
  XNR21 U2684 ( .A(n2820), .B(n2911), .Q(n3244) );
  OAI221 U2685 ( .A(n3245), .B(n2864), .C(n2965), .D(n3246), .Q(n1739) );
  XNR21 U2686 ( .A(n2821), .B(n2911), .Q(n3245) );
  OAI221 U2687 ( .A(n3246), .B(n2864), .C(n2965), .D(n3247), .Q(n1738) );
  XNR21 U2688 ( .A(n2822), .B(n2911), .Q(n3246) );
  OAI221 U2689 ( .A(n3247), .B(n2864), .C(n2965), .D(n3248), .Q(n1737) );
  XNR21 U2690 ( .A(n2823), .B(n2911), .Q(n3247) );
  OAI221 U2691 ( .A(n3248), .B(n2864), .C(n2965), .D(n3249), .Q(n1736) );
  XNR21 U2692 ( .A(n2824), .B(n2911), .Q(n3248) );
  OAI221 U2693 ( .A(n3249), .B(n2864), .C(n2965), .D(n3250), .Q(n1735) );
  XNR21 U2694 ( .A(n2825), .B(n2911), .Q(n3249) );
  OAI221 U2695 ( .A(n3250), .B(n2864), .C(n2965), .D(n3251), .Q(n1734) );
  XNR21 U2696 ( .A(n2826), .B(n2911), .Q(n3250) );
  OAI221 U2697 ( .A(n3251), .B(n2864), .C(n2965), .D(n3252), .Q(n1733) );
  XNR21 U2698 ( .A(n2827), .B(n2912), .Q(n3251) );
  OAI221 U2699 ( .A(n3252), .B(n2864), .C(n2965), .D(n3253), .Q(n1732) );
  XNR21 U2700 ( .A(n2828), .B(n2912), .Q(n3252) );
  OAI221 U2701 ( .A(n3253), .B(n2864), .C(n2965), .D(n3254), .Q(n1731) );
  XNR21 U2702 ( .A(n2829), .B(n2912), .Q(n3253) );
  OAI221 U2703 ( .A(n3254), .B(n2864), .C(n2965), .D(n3255), .Q(n1730) );
  XNR21 U2704 ( .A(n2830), .B(n2912), .Q(n3254) );
  OAI221 U2705 ( .A(n3255), .B(n2864), .C(n2965), .D(n3256), .Q(n1729) );
  XNR21 U2706 ( .A(n2831), .B(n2912), .Q(n3255) );
  OAI221 U2707 ( .A(n3256), .B(n2864), .C(n2965), .D(n3257), .Q(n1728) );
  XNR21 U2708 ( .A(n2832), .B(n2912), .Q(n3256) );
  OAI221 U2709 ( .A(n3257), .B(n2864), .C(n2965), .D(n3258), .Q(n1727) );
  XNR21 U2710 ( .A(n2833), .B(n2912), .Q(n3257) );
  OAI221 U2711 ( .A(n3258), .B(n2864), .C(n2965), .D(n3259), .Q(n1726) );
  XNR21 U2712 ( .A(n2834), .B(n2912), .Q(n3258) );
  OAI221 U2713 ( .A(n3259), .B(n2864), .C(n2965), .D(n3260), .Q(n1725) );
  XNR21 U2714 ( .A(n2835), .B(n2912), .Q(n3259) );
  OAI221 U2715 ( .A(n3260), .B(n2864), .C(n2965), .D(n3261), .Q(n1724) );
  XNR21 U2716 ( .A(n2836), .B(n2912), .Q(n3260) );
  OAI221 U2717 ( .A(n3261), .B(n2864), .C(n2965), .D(n3262), .Q(n1723) );
  XNR21 U2718 ( .A(n2837), .B(n2912), .Q(n3261) );
  OAI221 U2719 ( .A(n3262), .B(n2864), .C(n2965), .D(n3263), .Q(n1722) );
  XNR21 U2720 ( .A(n2838), .B(n2912), .Q(n3262) );
  OAI221 U2721 ( .A(n3263), .B(n2864), .C(n2965), .D(n3264), .Q(n1721) );
  XNR21 U2722 ( .A(n2839), .B(n2912), .Q(n3263) );
  OAI221 U2723 ( .A(n3264), .B(n2864), .C(n2965), .D(n3265), .Q(n1720) );
  XNR21 U2724 ( .A(n2840), .B(n2912), .Q(n3264) );
  OAI221 U2725 ( .A(n3265), .B(n2864), .C(n2965), .D(n3266), .Q(n1719) );
  XNR21 U2726 ( .A(n2841), .B(n2912), .Q(n3265) );
  OAI221 U2727 ( .A(n3266), .B(n2864), .C(n2965), .D(n3267), .Q(n1718) );
  XNR21 U2728 ( .A(n2842), .B(n2912), .Q(n3266) );
  OAI221 U2729 ( .A(n3267), .B(n2864), .C(n2965), .D(n3268), .Q(n1717) );
  XNR21 U2730 ( .A(n2843), .B(n2912), .Q(n3267) );
  OAI221 U2731 ( .A(n3268), .B(n2864), .C(n2965), .D(n3269), .Q(n1716) );
  XNR21 U2732 ( .A(n2844), .B(n2912), .Q(n3268) );
  OAI221 U2733 ( .A(n3269), .B(n2864), .C(n2965), .D(n3270), .Q(n1715) );
  XNR21 U2734 ( .A(n2845), .B(n2912), .Q(n3269) );
  OAI221 U2735 ( .A(n3270), .B(n2864), .C(n2965), .D(n3007), .Q(n1714) );
  XNR21 U2736 ( .A(n2847), .B(n2912), .Q(n3007) );
  XNR21 U2737 ( .A(n2846), .B(n2912), .Q(n3270) );
  AOI211 U2738 ( .A(n2864), .B(n2965), .C(n2741), .Q(n3271) );
  NOR22 U2739 ( .A(n2962), .B(n2849), .Q(n1712) );
  OAI221 U2740 ( .A(n3272), .B(n2865), .C(n2962), .D(n3273), .Q(n1711) );
  XNR21 U2741 ( .A(n2849), .B(n2916), .Q(n3272) );
  OAI221 U2742 ( .A(n3273), .B(n2865), .C(n2962), .D(n3274), .Q(n1710) );
  XNR21 U2743 ( .A(n2818), .B(n2914), .Q(n3273) );
  OAI221 U2744 ( .A(n3274), .B(n2865), .C(n2962), .D(n3275), .Q(n1709) );
  XNR21 U2745 ( .A(n2819), .B(n2914), .Q(n3274) );
  OAI221 U2746 ( .A(n3275), .B(n2865), .C(n2962), .D(n3276), .Q(n1708) );
  XNR21 U2747 ( .A(n2820), .B(n2914), .Q(n3275) );
  OAI221 U2748 ( .A(n3276), .B(n2865), .C(n2962), .D(n3277), .Q(n1707) );
  XNR21 U2749 ( .A(n2821), .B(n2914), .Q(n3276) );
  OAI221 U2750 ( .A(n3277), .B(n2865), .C(n2962), .D(n3278), .Q(n1706) );
  XNR21 U2751 ( .A(n2822), .B(n2914), .Q(n3277) );
  OAI221 U2752 ( .A(n3278), .B(n2866), .C(n2962), .D(n3279), .Q(n1705) );
  XNR21 U2753 ( .A(n2823), .B(n2914), .Q(n3278) );
  OAI221 U2754 ( .A(n3279), .B(n2866), .C(n2962), .D(n3280), .Q(n1704) );
  XNR21 U2755 ( .A(n2824), .B(n2914), .Q(n3279) );
  OAI221 U2756 ( .A(n3280), .B(n2866), .C(n2962), .D(n3281), .Q(n1703) );
  XNR21 U2757 ( .A(n2825), .B(n2914), .Q(n3280) );
  OAI221 U2758 ( .A(n3281), .B(n2866), .C(n2962), .D(n3282), .Q(n1702) );
  XNR21 U2759 ( .A(n2826), .B(n2914), .Q(n3281) );
  OAI221 U2760 ( .A(n3282), .B(n2866), .C(n2962), .D(n3283), .Q(n1701) );
  XNR21 U2761 ( .A(n2827), .B(n2915), .Q(n3282) );
  OAI221 U2762 ( .A(n3283), .B(n2866), .C(n2962), .D(n3284), .Q(n1700) );
  XNR21 U2763 ( .A(n2828), .B(n2915), .Q(n3283) );
  OAI221 U2764 ( .A(n3284), .B(n2866), .C(n2962), .D(n3285), .Q(n1699) );
  XNR21 U2765 ( .A(n2829), .B(n2915), .Q(n3284) );
  OAI221 U2766 ( .A(n3285), .B(n2867), .C(n2962), .D(n3286), .Q(n1698) );
  XNR21 U2767 ( .A(n2830), .B(n2915), .Q(n3285) );
  OAI221 U2768 ( .A(n3286), .B(n2867), .C(n2962), .D(n3287), .Q(n1697) );
  XNR21 U2769 ( .A(n2831), .B(n2915), .Q(n3286) );
  OAI221 U2770 ( .A(n3287), .B(n2867), .C(n2962), .D(n3288), .Q(n1696) );
  XNR21 U2771 ( .A(n2832), .B(n2915), .Q(n3287) );
  OAI221 U2772 ( .A(n3288), .B(n2867), .C(n2962), .D(n3289), .Q(n1695) );
  XNR21 U2773 ( .A(n2833), .B(n2915), .Q(n3288) );
  OAI221 U2774 ( .A(n3289), .B(n2867), .C(n2962), .D(n3290), .Q(n1694) );
  XNR21 U2775 ( .A(n2834), .B(n2915), .Q(n3289) );
  OAI221 U2776 ( .A(n3290), .B(n2867), .C(n2962), .D(n3291), .Q(n1693) );
  XNR21 U2777 ( .A(n2835), .B(n2915), .Q(n3290) );
  OAI221 U2778 ( .A(n3291), .B(n2868), .C(n2962), .D(n3292), .Q(n1692) );
  XNR21 U2779 ( .A(n2836), .B(n2915), .Q(n3291) );
  OAI221 U2780 ( .A(n3292), .B(n2868), .C(n2962), .D(n3293), .Q(n1691) );
  XNR21 U2781 ( .A(n2837), .B(n2915), .Q(n3292) );
  OAI221 U2782 ( .A(n3293), .B(n2868), .C(n2962), .D(n3294), .Q(n1690) );
  XNR21 U2783 ( .A(n2838), .B(n2915), .Q(n3293) );
  OAI221 U2784 ( .A(n3294), .B(n2868), .C(n2962), .D(n3295), .Q(n1689) );
  XNR21 U2785 ( .A(n2839), .B(n2915), .Q(n3294) );
  OAI221 U2786 ( .A(n3295), .B(n2868), .C(n2962), .D(n3296), .Q(n1688) );
  XNR21 U2787 ( .A(n2840), .B(n2915), .Q(n3295) );
  OAI221 U2788 ( .A(n3296), .B(n2868), .C(n2962), .D(n3297), .Q(n1687) );
  XNR21 U2789 ( .A(n2841), .B(n2915), .Q(n3296) );
  OAI221 U2790 ( .A(n3297), .B(n2868), .C(n2962), .D(n3298), .Q(n1686) );
  XNR21 U2791 ( .A(n2842), .B(n2915), .Q(n3297) );
  OAI221 U2792 ( .A(n3298), .B(n2869), .C(n2962), .D(n3299), .Q(n1685) );
  XNR21 U2793 ( .A(n2843), .B(n2915), .Q(n3298) );
  OAI221 U2794 ( .A(n3299), .B(n2869), .C(n2962), .D(n3300), .Q(n1684) );
  XNR21 U2795 ( .A(n2844), .B(n2915), .Q(n3299) );
  OAI221 U2796 ( .A(n3300), .B(n2869), .C(n2962), .D(n3301), .Q(n1683) );
  XNR21 U2797 ( .A(n2845), .B(n2915), .Q(n3300) );
  OAI221 U2798 ( .A(n3301), .B(n2869), .C(n2962), .D(n3009), .Q(n1682) );
  XNR21 U2799 ( .A(n2847), .B(n2915), .Q(n3009) );
  XNR21 U2800 ( .A(n2846), .B(n2915), .Q(n3301) );
  AOI211 U2801 ( .A(n2869), .B(n2962), .C(n2742), .Q(n3302) );
  NOR22 U2802 ( .A(n2959), .B(n2849), .Q(n1680) );
  OAI221 U2803 ( .A(n3303), .B(n2870), .C(n2959), .D(n3304), .Q(n1679) );
  XNR21 U2804 ( .A(n2849), .B(n2919), .Q(n3303) );
  OAI221 U2805 ( .A(n3304), .B(n3012), .C(n2959), .D(n3305), .Q(n1678) );
  XNR21 U2806 ( .A(n2818), .B(n2917), .Q(n3304) );
  OAI221 U2807 ( .A(n3305), .B(n2870), .C(n2959), .D(n3306), .Q(n1677) );
  XNR21 U2808 ( .A(n2819), .B(n2917), .Q(n3305) );
  OAI221 U2809 ( .A(n3306), .B(n2870), .C(n2959), .D(n3307), .Q(n1676) );
  XNR21 U2810 ( .A(n2820), .B(n2917), .Q(n3306) );
  OAI221 U2811 ( .A(n3307), .B(n3012), .C(n2959), .D(n3308), .Q(n1675) );
  XNR21 U2812 ( .A(n2821), .B(n2917), .Q(n3307) );
  OAI221 U2813 ( .A(n3308), .B(n3012), .C(n2959), .D(n3309), .Q(n1674) );
  XNR21 U2814 ( .A(n2822), .B(n2917), .Q(n3308) );
  OAI221 U2815 ( .A(n3309), .B(n3012), .C(n2959), .D(n3310), .Q(n1673) );
  XNR21 U2816 ( .A(n2823), .B(n2917), .Q(n3309) );
  OAI221 U2817 ( .A(n3310), .B(n3012), .C(n2959), .D(n3311), .Q(n1672) );
  XNR21 U2818 ( .A(n2824), .B(n2917), .Q(n3310) );
  OAI221 U2819 ( .A(n3311), .B(n3012), .C(n2959), .D(n3312), .Q(n1671) );
  XNR21 U2820 ( .A(n2825), .B(n2917), .Q(n3311) );
  OAI221 U2821 ( .A(n3312), .B(n3012), .C(n2959), .D(n3313), .Q(n1670) );
  XNR21 U2822 ( .A(n2826), .B(n2917), .Q(n3312) );
  OAI221 U2823 ( .A(n3313), .B(n3012), .C(n2959), .D(n3314), .Q(n1669) );
  XNR21 U2824 ( .A(n2827), .B(n2918), .Q(n3313) );
  OAI221 U2825 ( .A(n3314), .B(n3012), .C(n2959), .D(n3315), .Q(n1668) );
  XNR21 U2826 ( .A(n2828), .B(n2918), .Q(n3314) );
  OAI221 U2827 ( .A(n3315), .B(n3012), .C(n2959), .D(n3316), .Q(n1667) );
  XNR21 U2828 ( .A(n2829), .B(n2918), .Q(n3315) );
  OAI221 U2829 ( .A(n3316), .B(n3012), .C(n2959), .D(n3317), .Q(n1666) );
  XNR21 U2830 ( .A(n2830), .B(n2918), .Q(n3316) );
  OAI221 U2831 ( .A(n3317), .B(n3012), .C(n2959), .D(n3318), .Q(n1665) );
  XNR21 U2832 ( .A(n2831), .B(n2918), .Q(n3317) );
  OAI221 U2833 ( .A(n3318), .B(n3012), .C(n2959), .D(n3319), .Q(n1664) );
  XNR21 U2834 ( .A(n2832), .B(n2918), .Q(n3318) );
  OAI221 U2835 ( .A(n3319), .B(n3012), .C(n2959), .D(n3320), .Q(n1663) );
  XNR21 U2836 ( .A(n2833), .B(n2918), .Q(n3319) );
  OAI221 U2837 ( .A(n3320), .B(n3012), .C(n2959), .D(n3321), .Q(n1662) );
  XNR21 U2838 ( .A(n2834), .B(n2918), .Q(n3320) );
  OAI221 U2839 ( .A(n3321), .B(n2870), .C(n2959), .D(n3322), .Q(n1661) );
  XNR21 U2840 ( .A(n2835), .B(n2918), .Q(n3321) );
  OAI221 U2841 ( .A(n3322), .B(n3012), .C(n2959), .D(n3323), .Q(n1660) );
  XNR21 U2842 ( .A(n2836), .B(n2918), .Q(n3322) );
  OAI221 U2843 ( .A(n3323), .B(n3012), .C(n2959), .D(n3324), .Q(n1659) );
  XNR21 U2844 ( .A(n2837), .B(n2918), .Q(n3323) );
  OAI221 U2845 ( .A(n3324), .B(n3012), .C(n2959), .D(n3325), .Q(n1658) );
  XNR21 U2846 ( .A(n2838), .B(n2918), .Q(n3324) );
  OAI221 U2847 ( .A(n3325), .B(n2870), .C(n2959), .D(n3326), .Q(n1657) );
  XNR21 U2848 ( .A(n2839), .B(n2918), .Q(n3325) );
  OAI221 U2849 ( .A(n3326), .B(n2870), .C(n2959), .D(n3327), .Q(n1656) );
  XNR21 U2850 ( .A(n2840), .B(n2918), .Q(n3326) );
  OAI221 U2851 ( .A(n3327), .B(n2870), .C(n2959), .D(n3328), .Q(n1655) );
  XNR21 U2852 ( .A(n2841), .B(n2918), .Q(n3327) );
  OAI221 U2853 ( .A(n3328), .B(n2870), .C(n2959), .D(n3329), .Q(n1654) );
  XNR21 U2854 ( .A(n2842), .B(n2918), .Q(n3328) );
  OAI221 U2855 ( .A(n3329), .B(n2870), .C(n2959), .D(n3330), .Q(n1653) );
  XNR21 U2856 ( .A(n2843), .B(n2918), .Q(n3329) );
  OAI221 U2857 ( .A(n3330), .B(n2870), .C(n2959), .D(n3331), .Q(n1652) );
  XNR21 U2858 ( .A(n2844), .B(n2918), .Q(n3330) );
  OAI221 U2859 ( .A(n3331), .B(n2870), .C(n2959), .D(n3332), .Q(n1651) );
  XNR21 U2860 ( .A(n2845), .B(n2918), .Q(n3331) );
  OAI221 U2861 ( .A(n3332), .B(n2870), .C(n2959), .D(n3011), .Q(n1650) );
  XNR21 U2862 ( .A(n2847), .B(n2918), .Q(n3011) );
  XNR21 U2863 ( .A(n2846), .B(n2918), .Q(n3332) );
  AOI211 U2864 ( .A(n2870), .B(n2959), .C(n2743), .Q(n3333) );
  NOR22 U2865 ( .A(n2956), .B(n2986), .Q(n1648) );
  OAI221 U2866 ( .A(n3334), .B(n2871), .C(n2956), .D(n3335), .Q(n1647) );
  XNR21 U2867 ( .A(n2849), .B(n2922), .Q(n3334) );
  OAI221 U2868 ( .A(n3335), .B(n2871), .C(n2956), .D(n3336), .Q(n1646) );
  XNR21 U2869 ( .A(n2818), .B(n2920), .Q(n3335) );
  OAI221 U2870 ( .A(n3336), .B(n2871), .C(n2956), .D(n3337), .Q(n1645) );
  XNR21 U2871 ( .A(n2819), .B(n2920), .Q(n3336) );
  OAI221 U2872 ( .A(n3337), .B(n2871), .C(n2956), .D(n3338), .Q(n1644) );
  XNR21 U2873 ( .A(n2820), .B(n2920), .Q(n3337) );
  OAI221 U2874 ( .A(n3338), .B(n2871), .C(n2956), .D(n3339), .Q(n1643) );
  XNR21 U2875 ( .A(n2821), .B(n2920), .Q(n3338) );
  OAI221 U2876 ( .A(n3339), .B(n2871), .C(n2956), .D(n3340), .Q(n1642) );
  XNR21 U2877 ( .A(n2822), .B(n2920), .Q(n3339) );
  OAI221 U2878 ( .A(n3340), .B(n2872), .C(n2956), .D(n3341), .Q(n1641) );
  XNR21 U2879 ( .A(n2823), .B(n2920), .Q(n3340) );
  OAI221 U2880 ( .A(n3341), .B(n2872), .C(n2956), .D(n3342), .Q(n1640) );
  XNR21 U2881 ( .A(n2824), .B(n2920), .Q(n3341) );
  OAI221 U2882 ( .A(n3342), .B(n2872), .C(n2956), .D(n3343), .Q(n1639) );
  XNR21 U2883 ( .A(n2825), .B(n2920), .Q(n3342) );
  OAI221 U2884 ( .A(n3343), .B(n2872), .C(n2956), .D(n3344), .Q(n1638) );
  XNR21 U2885 ( .A(n2826), .B(n2920), .Q(n3343) );
  OAI221 U2886 ( .A(n3344), .B(n2872), .C(n2956), .D(n3345), .Q(n1637) );
  XNR21 U2887 ( .A(n2827), .B(n2921), .Q(n3344) );
  OAI221 U2888 ( .A(n3345), .B(n2872), .C(n2956), .D(n3346), .Q(n1636) );
  XNR21 U2889 ( .A(n2828), .B(n2921), .Q(n3345) );
  OAI221 U2890 ( .A(n3346), .B(n2872), .C(n2956), .D(n3347), .Q(n1635) );
  XNR21 U2891 ( .A(n2829), .B(n2921), .Q(n3346) );
  OAI221 U2892 ( .A(n3347), .B(n2873), .C(n2956), .D(n3348), .Q(n1634) );
  XNR21 U2893 ( .A(n2830), .B(n2921), .Q(n3347) );
  OAI221 U2894 ( .A(n3348), .B(n2873), .C(n2956), .D(n3349), .Q(n1633) );
  XNR21 U2895 ( .A(n2831), .B(n2921), .Q(n3348) );
  OAI221 U2896 ( .A(n3349), .B(n2873), .C(n2956), .D(n3350), .Q(n1632) );
  XNR21 U2897 ( .A(n2832), .B(n2921), .Q(n3349) );
  OAI221 U2898 ( .A(n3350), .B(n2873), .C(n2956), .D(n3351), .Q(n1631) );
  XNR21 U2899 ( .A(n2833), .B(n2921), .Q(n3350) );
  OAI221 U2900 ( .A(n3351), .B(n2873), .C(n2956), .D(n3352), .Q(n1630) );
  XNR21 U2901 ( .A(n2834), .B(n2921), .Q(n3351) );
  OAI221 U2902 ( .A(n3352), .B(n2873), .C(n2956), .D(n3353), .Q(n1629) );
  XNR21 U2903 ( .A(n2835), .B(n2921), .Q(n3352) );
  OAI221 U2904 ( .A(n3353), .B(n2874), .C(n2956), .D(n3354), .Q(n1628) );
  XNR21 U2905 ( .A(n2836), .B(n2921), .Q(n3353) );
  OAI221 U2906 ( .A(n3354), .B(n2874), .C(n2956), .D(n3355), .Q(n1627) );
  XNR21 U2907 ( .A(n2837), .B(n2921), .Q(n3354) );
  OAI221 U2908 ( .A(n3355), .B(n2874), .C(n2956), .D(n3356), .Q(n1626) );
  XNR21 U2909 ( .A(n2838), .B(n2921), .Q(n3355) );
  OAI221 U2910 ( .A(n3356), .B(n2874), .C(n2956), .D(n3357), .Q(n1625) );
  XNR21 U2911 ( .A(n2839), .B(n2921), .Q(n3356) );
  OAI221 U2912 ( .A(n3357), .B(n2874), .C(n2956), .D(n3358), .Q(n1624) );
  XNR21 U2913 ( .A(n2840), .B(n2921), .Q(n3357) );
  OAI221 U2914 ( .A(n3358), .B(n2874), .C(n2956), .D(n3359), .Q(n1623) );
  XNR21 U2915 ( .A(n2841), .B(n2921), .Q(n3358) );
  OAI221 U2916 ( .A(n3359), .B(n2874), .C(n2956), .D(n3360), .Q(n1622) );
  XNR21 U2917 ( .A(n2842), .B(n2921), .Q(n3359) );
  OAI221 U2918 ( .A(n3360), .B(n2875), .C(n2956), .D(n3361), .Q(n1621) );
  XNR21 U2919 ( .A(n2843), .B(n2921), .Q(n3360) );
  OAI221 U2920 ( .A(n3361), .B(n2875), .C(n2956), .D(n3362), .Q(n1620) );
  XNR21 U2921 ( .A(n2844), .B(n2921), .Q(n3361) );
  OAI221 U2922 ( .A(n3362), .B(n2875), .C(n2956), .D(n3363), .Q(n1619) );
  XNR21 U2923 ( .A(n2845), .B(n2921), .Q(n3362) );
  OAI221 U2924 ( .A(n3363), .B(n2875), .C(n2956), .D(n3013), .Q(n1618) );
  XNR21 U2925 ( .A(n2847), .B(n2921), .Q(n3013) );
  XNR21 U2926 ( .A(n2846), .B(n2921), .Q(n3363) );
  AOI211 U2927 ( .A(n2875), .B(n2956), .C(n2744), .Q(n3364) );
  NOR22 U2928 ( .A(n2953), .B(n2849), .Q(n1616) );
  OAI221 U2929 ( .A(n3365), .B(n2876), .C(n2953), .D(n3366), .Q(n1615) );
  XNR21 U2930 ( .A(n2849), .B(n2924), .Q(n3365) );
  OAI221 U2931 ( .A(n3366), .B(n2876), .C(n2953), .D(n3367), .Q(n1614) );
  XNR21 U2932 ( .A(n2818), .B(n2923), .Q(n3366) );
  OAI221 U2933 ( .A(n3367), .B(n2876), .C(n2953), .D(n3368), .Q(n1613) );
  XNR21 U2934 ( .A(n2819), .B(n2923), .Q(n3367) );
  OAI221 U2935 ( .A(n3368), .B(n2876), .C(n2953), .D(n3369), .Q(n1612) );
  XNR21 U2936 ( .A(n2820), .B(n2923), .Q(n3368) );
  OAI221 U2937 ( .A(n3369), .B(n2876), .C(n2953), .D(n3370), .Q(n1611) );
  XNR21 U2938 ( .A(n2821), .B(n2923), .Q(n3369) );
  OAI221 U2939 ( .A(n3370), .B(n2876), .C(n2953), .D(n3371), .Q(n1610) );
  XNR21 U2940 ( .A(n2822), .B(n2923), .Q(n3370) );
  OAI221 U2941 ( .A(n3371), .B(n2877), .C(n2953), .D(n3372), .Q(n1609) );
  XNR21 U2942 ( .A(n2823), .B(n2923), .Q(n3371) );
  OAI221 U2943 ( .A(n3372), .B(n2877), .C(n2953), .D(n3373), .Q(n1608) );
  XNR21 U2944 ( .A(n2824), .B(n2923), .Q(n3372) );
  OAI221 U2945 ( .A(n3373), .B(n2877), .C(n2953), .D(n3374), .Q(n1607) );
  XNR21 U2946 ( .A(n2825), .B(n2923), .Q(n3373) );
  OAI221 U2947 ( .A(n3374), .B(n2877), .C(n2953), .D(n3375), .Q(n1606) );
  XNR21 U2948 ( .A(n2826), .B(n2923), .Q(n3374) );
  OAI221 U2949 ( .A(n3375), .B(n2877), .C(n2953), .D(n3376), .Q(n1605) );
  XNR21 U2950 ( .A(n2827), .B(n2923), .Q(n3375) );
  OAI221 U2951 ( .A(n3376), .B(n2877), .C(n2953), .D(n3377), .Q(n1604) );
  XNR21 U2952 ( .A(n2828), .B(n2923), .Q(n3376) );
  OAI221 U2953 ( .A(n3377), .B(n2877), .C(n2953), .D(n3378), .Q(n1603) );
  XNR21 U2954 ( .A(n2829), .B(n2923), .Q(n3377) );
  OAI221 U2955 ( .A(n3378), .B(n2878), .C(n2953), .D(n3379), .Q(n1602) );
  XNR21 U2956 ( .A(n2830), .B(n2923), .Q(n3378) );
  OAI221 U2957 ( .A(n3379), .B(n2878), .C(n2953), .D(n3380), .Q(n1601) );
  XNR21 U2958 ( .A(n2831), .B(n2923), .Q(n3379) );
  OAI221 U2959 ( .A(n3380), .B(n2878), .C(n2953), .D(n3381), .Q(n1600) );
  XNR21 U2960 ( .A(n2832), .B(n2923), .Q(n3380) );
  OAI221 U2961 ( .A(n3381), .B(n2878), .C(n2953), .D(n3382), .Q(n1599) );
  XNR21 U2962 ( .A(n2833), .B(n2923), .Q(n3381) );
  OAI221 U2963 ( .A(n3382), .B(n2878), .C(n2953), .D(n3383), .Q(n1598) );
  XNR21 U2964 ( .A(n2834), .B(n2923), .Q(n3382) );
  OAI221 U2965 ( .A(n3383), .B(n2878), .C(n2953), .D(n3384), .Q(n1597) );
  XNR21 U2966 ( .A(n2835), .B(n2923), .Q(n3383) );
  OAI221 U2967 ( .A(n3384), .B(n2879), .C(n2953), .D(n3385), .Q(n1596) );
  XNR21 U2968 ( .A(n2836), .B(n2923), .Q(n3384) );
  OAI221 U2969 ( .A(n3385), .B(n2879), .C(n2953), .D(n3386), .Q(n1595) );
  XNR21 U2970 ( .A(n2837), .B(n2923), .Q(n3385) );
  OAI221 U2971 ( .A(n3386), .B(n2879), .C(n2953), .D(n3387), .Q(n1594) );
  XNR21 U2972 ( .A(n2838), .B(n2923), .Q(n3386) );
  OAI221 U2973 ( .A(n3387), .B(n2879), .C(n2953), .D(n3388), .Q(n1593) );
  XNR21 U2974 ( .A(n2839), .B(n2923), .Q(n3387) );
  OAI221 U2975 ( .A(n3388), .B(n2879), .C(n2953), .D(n3389), .Q(n1592) );
  XNR21 U2976 ( .A(n2840), .B(n2923), .Q(n3388) );
  OAI221 U2977 ( .A(n3389), .B(n2879), .C(n2953), .D(n3390), .Q(n1591) );
  XNR21 U2978 ( .A(n2841), .B(n2923), .Q(n3389) );
  OAI221 U2979 ( .A(n3390), .B(n2879), .C(n2953), .D(n3391), .Q(n1590) );
  XNR21 U2980 ( .A(n2842), .B(n2923), .Q(n3390) );
  OAI221 U2981 ( .A(n3391), .B(n2880), .C(n2953), .D(n3392), .Q(n1589) );
  XNR21 U2982 ( .A(n2843), .B(n2923), .Q(n3391) );
  OAI221 U2983 ( .A(n3392), .B(n2880), .C(n2953), .D(n3393), .Q(n1588) );
  XNR21 U2984 ( .A(n2844), .B(a[23]), .Q(n3392) );
  OAI221 U2985 ( .A(n3393), .B(n2880), .C(n2953), .D(n3394), .Q(n1587) );
  XNR21 U2986 ( .A(n2845), .B(a[23]), .Q(n3393) );
  OAI221 U2987 ( .A(n3394), .B(n2880), .C(n2953), .D(n3015), .Q(n1586) );
  XNR21 U2988 ( .A(n2847), .B(a[23]), .Q(n3015) );
  XNR21 U2989 ( .A(n2846), .B(a[23]), .Q(n3394) );
  AOI211 U2990 ( .A(n2880), .B(n2953), .C(n2745), .Q(n3395) );
  NOR22 U2991 ( .A(n2950), .B(n2986), .Q(n1584) );
  OAI221 U2992 ( .A(n3396), .B(n2881), .C(n2950), .D(n3397), .Q(n1583) );
  XNR21 U2993 ( .A(n2849), .B(n2927), .Q(n3396) );
  OAI221 U2994 ( .A(n3397), .B(n2881), .C(n2950), .D(n3398), .Q(n1582) );
  XNR21 U2995 ( .A(n2818), .B(n2925), .Q(n3397) );
  OAI221 U2996 ( .A(n3398), .B(n2881), .C(n2950), .D(n3399), .Q(n1581) );
  XNR21 U2997 ( .A(n2819), .B(n2925), .Q(n3398) );
  OAI221 U2998 ( .A(n3399), .B(n2881), .C(n2950), .D(n3400), .Q(n1580) );
  XNR21 U2999 ( .A(n2820), .B(n2925), .Q(n3399) );
  OAI221 U3000 ( .A(n3400), .B(n2881), .C(n2950), .D(n3401), .Q(n1579) );
  XNR21 U3001 ( .A(n2821), .B(n2925), .Q(n3400) );
  OAI221 U3002 ( .A(n3401), .B(n2881), .C(n2950), .D(n3402), .Q(n1578) );
  XNR21 U3003 ( .A(n2822), .B(n2925), .Q(n3401) );
  OAI221 U3004 ( .A(n3402), .B(n2882), .C(n2950), .D(n3403), .Q(n1577) );
  XNR21 U3005 ( .A(n2823), .B(n2925), .Q(n3402) );
  OAI221 U3006 ( .A(n3403), .B(n2882), .C(n2950), .D(n3404), .Q(n1576) );
  XNR21 U3007 ( .A(n2824), .B(n2925), .Q(n3403) );
  OAI221 U3008 ( .A(n3404), .B(n2882), .C(n2950), .D(n3405), .Q(n1575) );
  XNR21 U3009 ( .A(n2825), .B(n2925), .Q(n3404) );
  OAI221 U3010 ( .A(n3405), .B(n2882), .C(n2950), .D(n3406), .Q(n1574) );
  XNR21 U3011 ( .A(n2826), .B(n2925), .Q(n3405) );
  OAI221 U3012 ( .A(n3406), .B(n2882), .C(n2950), .D(n3407), .Q(n1573) );
  XNR21 U3013 ( .A(n2827), .B(n2926), .Q(n3406) );
  OAI221 U3014 ( .A(n3407), .B(n2882), .C(n2950), .D(n3408), .Q(n1572) );
  XNR21 U3015 ( .A(n2828), .B(n2926), .Q(n3407) );
  OAI221 U3016 ( .A(n3408), .B(n2882), .C(n2950), .D(n3409), .Q(n1571) );
  XNR21 U3017 ( .A(n2829), .B(n2926), .Q(n3408) );
  OAI221 U3018 ( .A(n3409), .B(n2883), .C(n2950), .D(n3410), .Q(n1570) );
  XNR21 U3019 ( .A(n2830), .B(n2926), .Q(n3409) );
  OAI221 U3020 ( .A(n3410), .B(n2883), .C(n2950), .D(n3411), .Q(n1569) );
  XNR21 U3021 ( .A(n2831), .B(n2926), .Q(n3410) );
  OAI221 U3022 ( .A(n3411), .B(n2883), .C(n2950), .D(n3412), .Q(n1568) );
  XNR21 U3023 ( .A(n2832), .B(n2926), .Q(n3411) );
  OAI221 U3024 ( .A(n3412), .B(n2883), .C(n2950), .D(n3413), .Q(n1567) );
  XNR21 U3025 ( .A(n2833), .B(n2926), .Q(n3412) );
  OAI221 U3026 ( .A(n3413), .B(n2883), .C(n2950), .D(n3414), .Q(n1566) );
  XNR21 U3027 ( .A(n2834), .B(n2926), .Q(n3413) );
  OAI221 U3028 ( .A(n3414), .B(n2883), .C(n2950), .D(n3415), .Q(n1565) );
  XNR21 U3029 ( .A(n2835), .B(n2926), .Q(n3414) );
  OAI221 U3030 ( .A(n3415), .B(n2884), .C(n2950), .D(n3416), .Q(n1564) );
  XNR21 U3031 ( .A(n2836), .B(n2926), .Q(n3415) );
  OAI221 U3032 ( .A(n3416), .B(n2884), .C(n2950), .D(n3417), .Q(n1563) );
  XNR21 U3033 ( .A(n2837), .B(n2926), .Q(n3416) );
  OAI221 U3034 ( .A(n3417), .B(n2884), .C(n2950), .D(n3418), .Q(n1562) );
  XNR21 U3035 ( .A(n2838), .B(n2926), .Q(n3417) );
  OAI221 U3036 ( .A(n3418), .B(n2884), .C(n2950), .D(n3419), .Q(n1561) );
  XNR21 U3037 ( .A(n2839), .B(n2926), .Q(n3418) );
  OAI221 U3038 ( .A(n3419), .B(n2884), .C(n2950), .D(n3420), .Q(n1560) );
  XNR21 U3039 ( .A(n2840), .B(n2926), .Q(n3419) );
  OAI221 U3040 ( .A(n3420), .B(n2884), .C(n2950), .D(n3421), .Q(n1559) );
  XNR21 U3041 ( .A(n2841), .B(n2926), .Q(n3420) );
  OAI221 U3042 ( .A(n3421), .B(n2884), .C(n2950), .D(n3422), .Q(n1558) );
  XNR21 U3043 ( .A(n2842), .B(n2926), .Q(n3421) );
  OAI221 U3044 ( .A(n3422), .B(n2885), .C(n2950), .D(n3423), .Q(n1557) );
  XNR21 U3045 ( .A(n2843), .B(n2926), .Q(n3422) );
  OAI221 U3046 ( .A(n3423), .B(n2885), .C(n2950), .D(n3424), .Q(n1556) );
  XNR21 U3047 ( .A(n2844), .B(n2926), .Q(n3423) );
  OAI221 U3048 ( .A(n3424), .B(n2885), .C(n2950), .D(n3425), .Q(n1555) );
  XNR21 U3049 ( .A(n2845), .B(n2926), .Q(n3424) );
  OAI221 U3050 ( .A(n3425), .B(n2885), .C(n2950), .D(n3017), .Q(n1554) );
  XNR21 U3051 ( .A(n2847), .B(n2926), .Q(n3017) );
  XNR21 U3052 ( .A(n2846), .B(n2926), .Q(n3425) );
  AOI211 U3053 ( .A(n2885), .B(n2950), .C(n2746), .Q(n3426) );
  NOR22 U3054 ( .A(n2947), .B(n2986), .Q(n1552) );
  OAI221 U3055 ( .A(n3427), .B(n3020), .C(n2947), .D(n3428), .Q(n1551) );
  XNR21 U3056 ( .A(n2849), .B(n2930), .Q(n3427) );
  OAI221 U3057 ( .A(n3428), .B(n3020), .C(n2947), .D(n3429), .Q(n1550) );
  XNR21 U3058 ( .A(n2818), .B(n2928), .Q(n3428) );
  OAI221 U3059 ( .A(n3429), .B(n2886), .C(n2947), .D(n3430), .Q(n1549) );
  XNR21 U3060 ( .A(n2819), .B(n2928), .Q(n3429) );
  OAI221 U3061 ( .A(n3430), .B(n2889), .C(n2947), .D(n3431), .Q(n1548) );
  XNR21 U3062 ( .A(n2820), .B(n2928), .Q(n3430) );
  OAI221 U3063 ( .A(n3431), .B(n2888), .C(n2947), .D(n3432), .Q(n1547) );
  XNR21 U3064 ( .A(n2821), .B(n2928), .Q(n3431) );
  OAI221 U3065 ( .A(n3432), .B(n2887), .C(n2947), .D(n3433), .Q(n1546) );
  XNR21 U3066 ( .A(n2822), .B(n2928), .Q(n3432) );
  OAI221 U3067 ( .A(n3433), .B(n2886), .C(n2947), .D(n3434), .Q(n1545) );
  XNR21 U3068 ( .A(n2823), .B(n2928), .Q(n3433) );
  OAI221 U3069 ( .A(n3434), .B(n2886), .C(n2947), .D(n3435), .Q(n1544) );
  XNR21 U3070 ( .A(n2824), .B(n2928), .Q(n3434) );
  OAI221 U3071 ( .A(n3435), .B(n2886), .C(n2947), .D(n3436), .Q(n1543) );
  XNR21 U3072 ( .A(n2825), .B(n2928), .Q(n3435) );
  OAI221 U3073 ( .A(n3436), .B(n2886), .C(n2947), .D(n3437), .Q(n1542) );
  XNR21 U3074 ( .A(n2826), .B(n2928), .Q(n3436) );
  OAI221 U3075 ( .A(n3437), .B(n2886), .C(n2947), .D(n3438), .Q(n1541) );
  XNR21 U3076 ( .A(n2827), .B(n2929), .Q(n3437) );
  OAI221 U3077 ( .A(n3438), .B(n2886), .C(n2947), .D(n3439), .Q(n1540) );
  XNR21 U3078 ( .A(n2828), .B(n2929), .Q(n3438) );
  OAI221 U3079 ( .A(n3439), .B(n2886), .C(n2947), .D(n3440), .Q(n1539) );
  XNR21 U3080 ( .A(n2829), .B(n2929), .Q(n3439) );
  OAI221 U3081 ( .A(n3440), .B(n2887), .C(n2947), .D(n3441), .Q(n1538) );
  XNR21 U3082 ( .A(n2830), .B(n2929), .Q(n3440) );
  OAI221 U3083 ( .A(n3441), .B(n2887), .C(n2947), .D(n3442), .Q(n1537) );
  XNR21 U3084 ( .A(n2831), .B(n2929), .Q(n3441) );
  OAI221 U3085 ( .A(n3442), .B(n2887), .C(n2947), .D(n3443), .Q(n1536) );
  XNR21 U3086 ( .A(n2832), .B(n2929), .Q(n3442) );
  OAI221 U3087 ( .A(n3443), .B(n2887), .C(n2947), .D(n3444), .Q(n1535) );
  XNR21 U3088 ( .A(n2833), .B(n2929), .Q(n3443) );
  OAI221 U3089 ( .A(n3444), .B(n2887), .C(n2947), .D(n3445), .Q(n1534) );
  XNR21 U3090 ( .A(n2834), .B(n2929), .Q(n3444) );
  OAI221 U3091 ( .A(n3445), .B(n2887), .C(n2947), .D(n3446), .Q(n1533) );
  XNR21 U3092 ( .A(n2835), .B(n2929), .Q(n3445) );
  OAI221 U3093 ( .A(n3446), .B(n2888), .C(n2947), .D(n3447), .Q(n1532) );
  XNR21 U3094 ( .A(n2836), .B(n2929), .Q(n3446) );
  OAI221 U3095 ( .A(n3447), .B(n2888), .C(n2947), .D(n3448), .Q(n1531) );
  XNR21 U3096 ( .A(n2837), .B(n2929), .Q(n3447) );
  OAI221 U3097 ( .A(n3448), .B(n2888), .C(n2947), .D(n3449), .Q(n1530) );
  XNR21 U3098 ( .A(n2838), .B(n2929), .Q(n3448) );
  OAI221 U3099 ( .A(n3449), .B(n2888), .C(n2947), .D(n3450), .Q(n1529) );
  XNR21 U3100 ( .A(n2839), .B(n2929), .Q(n3449) );
  OAI221 U3101 ( .A(n3450), .B(n2888), .C(n2947), .D(n3451), .Q(n1528) );
  XNR21 U3102 ( .A(n2840), .B(n2929), .Q(n3450) );
  OAI221 U3103 ( .A(n3451), .B(n2888), .C(n2947), .D(n3452), .Q(n1527) );
  XNR21 U3104 ( .A(n2841), .B(n2929), .Q(n3451) );
  OAI221 U3105 ( .A(n3452), .B(n2888), .C(n2947), .D(n3453), .Q(n1526) );
  XNR21 U3106 ( .A(n2842), .B(n2929), .Q(n3452) );
  OAI221 U3107 ( .A(n3453), .B(n2889), .C(n2947), .D(n3454), .Q(n1525) );
  XNR21 U3108 ( .A(n2843), .B(n2929), .Q(n3453) );
  OAI221 U3109 ( .A(n3454), .B(n2889), .C(n2947), .D(n3455), .Q(n1524) );
  XNR21 U3110 ( .A(n2844), .B(n2929), .Q(n3454) );
  OAI221 U3111 ( .A(n3455), .B(n2889), .C(n2947), .D(n3456), .Q(n1523) );
  XNR21 U3112 ( .A(n2845), .B(n2929), .Q(n3455) );
  OAI221 U3113 ( .A(n3456), .B(n2889), .C(n2947), .D(n3019), .Q(n1522) );
  XNR21 U3114 ( .A(n2847), .B(n2929), .Q(n3019) );
  XNR21 U3115 ( .A(n2846), .B(n2929), .Q(n3456) );
  AOI211 U3116 ( .A(n2889), .B(n2947), .C(n2747), .Q(n3457) );
  NOR22 U3117 ( .A(n2944), .B(n2986), .Q(n1520) );
  OAI221 U3118 ( .A(n3458), .B(n2851), .C(n2944), .D(n3459), .Q(n1519) );
  XNR21 U3119 ( .A(n2849), .B(n2933), .Q(n3458) );
  OAI221 U3120 ( .A(n3459), .B(n2851), .C(n2944), .D(n3460), .Q(n1518) );
  XNR21 U3121 ( .A(n2818), .B(n2931), .Q(n3459) );
  OAI221 U3122 ( .A(n3460), .B(n2851), .C(n2944), .D(n2990), .Q(n1517) );
  XNR21 U3123 ( .A(n2820), .B(n2931), .Q(n2990) );
  XNR21 U3124 ( .A(n2819), .B(n2931), .Q(n3460) );
  OAI221 U3125 ( .A(n2992), .B(n2851), .C(n2944), .D(n3461), .Q(n1515) );
  XNR21 U3126 ( .A(n2821), .B(n2931), .Q(n2992) );
  OAI221 U3127 ( .A(n3461), .B(n2851), .C(n2944), .D(n3462), .Q(n1514) );
  XNR21 U3128 ( .A(n2822), .B(n2931), .Q(n3461) );
  OAI221 U3129 ( .A(n3462), .B(n2852), .C(n2944), .D(n3463), .Q(n1513) );
  XNR21 U3130 ( .A(n2823), .B(n2931), .Q(n3462) );
  OAI221 U3131 ( .A(n3463), .B(n2852), .C(n2944), .D(n3464), .Q(n1512) );
  XNR21 U3132 ( .A(n2824), .B(n2931), .Q(n3463) );
  OAI221 U3133 ( .A(n3464), .B(n2852), .C(n2944), .D(n3465), .Q(n1511) );
  XNR21 U3134 ( .A(n2825), .B(n2931), .Q(n3464) );
  OAI221 U3135 ( .A(n3465), .B(n2852), .C(n2944), .D(n3466), .Q(n1510) );
  XNR21 U3136 ( .A(n2826), .B(n2931), .Q(n3465) );
  OAI221 U3137 ( .A(n3466), .B(n2852), .C(n2944), .D(n3467), .Q(n1509) );
  XNR21 U3138 ( .A(n2827), .B(n2932), .Q(n3466) );
  OAI221 U3139 ( .A(n3467), .B(n2852), .C(n2944), .D(n3468), .Q(n1508) );
  XNR21 U3140 ( .A(n2828), .B(n2932), .Q(n3467) );
  OAI221 U3141 ( .A(n3468), .B(n2852), .C(n2944), .D(n3469), .Q(n1507) );
  XNR21 U3142 ( .A(n2829), .B(n2932), .Q(n3468) );
  OAI221 U3143 ( .A(n3469), .B(n2853), .C(n2944), .D(n3470), .Q(n1506) );
  XNR21 U3144 ( .A(n2830), .B(n2932), .Q(n3469) );
  OAI221 U3145 ( .A(n3470), .B(n2853), .C(n2944), .D(n3471), .Q(n1505) );
  XNR21 U3146 ( .A(n2831), .B(n2932), .Q(n3470) );
  OAI221 U3147 ( .A(n3471), .B(n2853), .C(n2944), .D(n3472), .Q(n1504) );
  XNR21 U3148 ( .A(n2832), .B(n2932), .Q(n3471) );
  OAI221 U3149 ( .A(n3472), .B(n2853), .C(n2944), .D(n3473), .Q(n1503) );
  XNR21 U3150 ( .A(n2833), .B(n2932), .Q(n3472) );
  OAI221 U3151 ( .A(n3473), .B(n2853), .C(n2944), .D(n3474), .Q(n1502) );
  XNR21 U3152 ( .A(n2834), .B(n2932), .Q(n3473) );
  OAI221 U3153 ( .A(n3474), .B(n2853), .C(n2944), .D(n3475), .Q(n1501) );
  XNR21 U3154 ( .A(n2835), .B(n2932), .Q(n3474) );
  OAI221 U3155 ( .A(n3475), .B(n2854), .C(n2944), .D(n3476), .Q(n1500) );
  XNR21 U3156 ( .A(n2836), .B(n2932), .Q(n3475) );
  OAI221 U3157 ( .A(n3476), .B(n2854), .C(n2944), .D(n3477), .Q(n1499) );
  XNR21 U3158 ( .A(n2837), .B(n2932), .Q(n3476) );
  OAI221 U3159 ( .A(n3477), .B(n2854), .C(n2944), .D(n3478), .Q(n1498) );
  XNR21 U3160 ( .A(n2838), .B(n2932), .Q(n3477) );
  OAI221 U3161 ( .A(n3478), .B(n2854), .C(n2944), .D(n3479), .Q(n1497) );
  XNR21 U3162 ( .A(n2839), .B(n2932), .Q(n3478) );
  OAI221 U3163 ( .A(n3479), .B(n2854), .C(n2944), .D(n3480), .Q(n1496) );
  XNR21 U3164 ( .A(n2840), .B(n2932), .Q(n3479) );
  OAI221 U3165 ( .A(n3480), .B(n2854), .C(n2944), .D(n3481), .Q(n1495) );
  XNR21 U3166 ( .A(n2841), .B(n2932), .Q(n3480) );
  OAI221 U3167 ( .A(n3481), .B(n2854), .C(n2944), .D(n3482), .Q(n1494) );
  XNR21 U3168 ( .A(n2842), .B(n2932), .Q(n3481) );
  OAI221 U3169 ( .A(n3482), .B(n2855), .C(n2944), .D(n3483), .Q(n1493) );
  XNR21 U3170 ( .A(n2843), .B(n2932), .Q(n3482) );
  OAI221 U3171 ( .A(n3483), .B(n2855), .C(n2944), .D(n3484), .Q(n1492) );
  XNR21 U3172 ( .A(n2844), .B(n2932), .Q(n3483) );
  OAI221 U3173 ( .A(n3484), .B(n2855), .C(n2944), .D(n3485), .Q(n1491) );
  XNR21 U3174 ( .A(n2845), .B(n2932), .Q(n3484) );
  OAI221 U3175 ( .A(n3485), .B(n2855), .C(n2944), .D(n3021), .Q(n1490) );
  XNR21 U3176 ( .A(n2847), .B(n2932), .Q(n3021) );
  XNR21 U3177 ( .A(n2846), .B(n2932), .Q(n3485) );
  AOI211 U3178 ( .A(n2855), .B(n2944), .C(n2748), .Q(n3486) );
  NOR22 U3179 ( .A(n2940), .B(n2986), .Q(n1488) );
  OAI221 U3180 ( .A(n3487), .B(n3023), .C(n2940), .D(n3488), .Q(n1487) );
  XNR21 U3181 ( .A(n2849), .B(n2936), .Q(n3487) );
  OAI221 U3182 ( .A(n3488), .B(n3023), .C(n2940), .D(n3489), .Q(n1486) );
  XNR21 U3183 ( .A(n2818), .B(n2934), .Q(n3488) );
  OAI221 U3184 ( .A(n3489), .B(n2890), .C(n2940), .D(n3490), .Q(n1485) );
  XNR21 U3185 ( .A(n2819), .B(n2934), .Q(n3489) );
  OAI221 U3186 ( .A(n3490), .B(n2890), .C(n2940), .D(n3491), .Q(n1484) );
  XNR21 U3187 ( .A(n2820), .B(n2934), .Q(n3490) );
  OAI221 U3188 ( .A(n3491), .B(n2890), .C(n2940), .D(n3492), .Q(n1483) );
  XNR21 U3189 ( .A(n2821), .B(n2934), .Q(n3491) );
  OAI221 U3190 ( .A(n3492), .B(n2890), .C(n2940), .D(n3493), .Q(n1482) );
  XNR21 U3191 ( .A(n2822), .B(n2934), .Q(n3492) );
  OAI221 U3192 ( .A(n3493), .B(n2890), .C(n2940), .D(n3494), .Q(n1481) );
  XNR21 U3193 ( .A(n2823), .B(n2934), .Q(n3493) );
  OAI221 U3194 ( .A(n3494), .B(n2890), .C(n2940), .D(n3495), .Q(n1480) );
  XNR21 U3195 ( .A(n2824), .B(n2934), .Q(n3494) );
  OAI221 U3196 ( .A(n3495), .B(n2890), .C(n2940), .D(n3496), .Q(n1479) );
  XNR21 U3197 ( .A(n2825), .B(n2934), .Q(n3495) );
  OAI221 U3198 ( .A(n3496), .B(n2890), .C(n2940), .D(n3497), .Q(n1478) );
  XNR21 U3199 ( .A(n2826), .B(n2934), .Q(n3496) );
  OAI221 U3200 ( .A(n3497), .B(n2890), .C(n2940), .D(n3498), .Q(n1477) );
  XNR21 U3201 ( .A(n2827), .B(n2935), .Q(n3497) );
  OAI221 U3202 ( .A(n3498), .B(n2890), .C(n2940), .D(n3499), .Q(n1476) );
  XNR21 U3203 ( .A(n2828), .B(n2935), .Q(n3498) );
  OAI221 U3204 ( .A(n3499), .B(n2890), .C(n2940), .D(n3500), .Q(n1475) );
  XNR21 U3205 ( .A(n2829), .B(n2935), .Q(n3499) );
  OAI221 U3206 ( .A(n3500), .B(n2890), .C(n2940), .D(n3501), .Q(n1474) );
  XNR21 U3207 ( .A(n2830), .B(n2935), .Q(n3500) );
  OAI221 U3208 ( .A(n3501), .B(n2890), .C(n2940), .D(n3502), .Q(n1473) );
  XNR21 U3209 ( .A(n2831), .B(n2935), .Q(n3501) );
  OAI221 U3210 ( .A(n3502), .B(n2890), .C(n2940), .D(n3503), .Q(n1472) );
  XNR21 U3211 ( .A(n2832), .B(n2935), .Q(n3502) );
  OAI221 U3212 ( .A(n3503), .B(n2890), .C(n2940), .D(n3504), .Q(n1471) );
  XNR21 U3213 ( .A(n2833), .B(n2935), .Q(n3503) );
  OAI221 U3214 ( .A(n3504), .B(n2890), .C(n2940), .D(n3505), .Q(n1470) );
  XNR21 U3215 ( .A(n2834), .B(n2935), .Q(n3504) );
  OAI221 U3216 ( .A(n3505), .B(n2890), .C(n2940), .D(n3506), .Q(n1469) );
  XNR21 U3217 ( .A(n2835), .B(n2935), .Q(n3505) );
  OAI221 U3218 ( .A(n3506), .B(n2890), .C(n2940), .D(n3507), .Q(n1468) );
  XNR21 U3219 ( .A(n2836), .B(n2935), .Q(n3506) );
  XNR21 U3220 ( .A(n2837), .B(n2935), .Q(n3507) );
  XNR21 U3221 ( .A(n2838), .B(n2935), .Q(n3508) );
  XNR21 U3222 ( .A(n2839), .B(n2935), .Q(n3509) );
  XNR21 U3223 ( .A(n2840), .B(n2935), .Q(n3510) );
  XNR21 U3224 ( .A(n2841), .B(n2935), .Q(n3511) );
  XNR21 U3225 ( .A(n2842), .B(n2935), .Q(n3512) );
  OAI221 U3226 ( .A(n3513), .B(n2890), .C(n2940), .D(n3514), .Q(n1461) );
  XNR21 U3227 ( .A(n2843), .B(n2935), .Q(n3513) );
  OAI221 U3228 ( .A(n3514), .B(n2890), .C(n2940), .D(n3515), .Q(n1460) );
  XNR21 U3229 ( .A(n2844), .B(n2935), .Q(n3514) );
  OAI221 U3230 ( .A(n3515), .B(n2890), .C(n2940), .D(n3516), .Q(n1459) );
  XNR21 U3231 ( .A(n2845), .B(n2935), .Q(n3515) );
  OAI221 U3232 ( .A(n3516), .B(n2890), .C(n2940), .D(n3022), .Q(n1458) );
  XNR21 U3233 ( .A(n2847), .B(n2935), .Q(n3022) );
  XNR21 U3234 ( .A(n2846), .B(n2935), .Q(n3516) );
  AOI211 U3235 ( .A(n2890), .B(n2940), .C(n2749), .Q(n3517) );
  OAI211 U3236 ( .A(b[0]), .B(n2894), .C(n3024), .Q(n1456) );
  OAI221 U3237 ( .A(n2897), .B(n2997), .C(n2897), .D(n3518), .Q(n1455) );
  NAND22 U3238 ( .A(n3519), .B(n2850), .Q(n3518) );
  XNR21 U3239 ( .A(a[4]), .B(n2900), .Q(n3523) );
  OAI221 U3240 ( .A(n2903), .B(n3001), .C(n2903), .D(n3524), .Q(n1453) );
  NAND22 U3241 ( .A(n3525), .B(n2849), .Q(n3524) );
  XNR21 U3242 ( .A(a[6]), .B(n2903), .Q(n3526) );
  OAI221 U3243 ( .A(n2906), .B(n3003), .C(n2906), .D(n3527), .Q(n1452) );
  NAND22 U3244 ( .A(n3528), .B(n2849), .Q(n3527) );
  NAND22 U3245 ( .A(n2974), .B(n3529), .Q(n3003) );
  XNR21 U3246 ( .A(a[8]), .B(n2906), .Q(n3529) );
  OAI221 U3247 ( .A(n2908), .B(n3005), .C(n2908), .D(n3530), .Q(n1451) );
  NAND22 U3248 ( .A(n3531), .B(n2849), .Q(n3530) );
  XNR21 U3249 ( .A(a[10]), .B(n2908), .Q(n3532) );
  XNR21 U3250 ( .A(n2906), .B(a[10]), .Q(n3531) );
  OAI221 U3251 ( .A(n2910), .B(n2994), .C(n2910), .D(n3533), .Q(n1450) );
  NAND22 U3252 ( .A(n3534), .B(n2849), .Q(n3533) );
  XNR21 U3253 ( .A(a[12]), .B(n2910), .Q(n3535) );
  XNR21 U3254 ( .A(a[12]), .B(n2908), .Q(n3534) );
  OAI221 U3255 ( .A(n2913), .B(n3008), .C(n2913), .D(n3536), .Q(n1449) );
  NAND22 U3256 ( .A(n3537), .B(n2849), .Q(n3536) );
  NAND22 U3257 ( .A(n2965), .B(n3538), .Q(n3008) );
  XNR21 U3258 ( .A(a[14]), .B(n2913), .Q(n3538) );
  XNR21 U3259 ( .A(a[14]), .B(n2910), .Q(n3537) );
  OAI221 U3260 ( .A(n2916), .B(n2865), .C(n2916), .D(n3539), .Q(n1448) );
  NAND22 U3261 ( .A(n3540), .B(n2850), .Q(n3539) );
  NAND22 U3262 ( .A(n2962), .B(n3541), .Q(n3010) );
  XNR21 U3263 ( .A(a[16]), .B(n2916), .Q(n3541) );
  XNR21 U3264 ( .A(a[16]), .B(n2913), .Q(n3540) );
  OAI221 U3265 ( .A(n2919), .B(n3012), .C(n2919), .D(n3542), .Q(n1447) );
  NAND22 U3266 ( .A(n3543), .B(n2850), .Q(n3542) );
  XNR21 U3267 ( .A(a[18]), .B(n2919), .Q(n3544) );
  XNR21 U3268 ( .A(a[18]), .B(n2916), .Q(n3543) );
  OAI221 U3269 ( .A(n2922), .B(n2871), .C(n2922), .D(n3545), .Q(n1446) );
  NAND22 U3270 ( .A(n3546), .B(n2850), .Q(n3545) );
  NAND22 U3271 ( .A(n2956), .B(n3547), .Q(n3014) );
  XNR21 U3272 ( .A(a[20]), .B(n2922), .Q(n3547) );
  XNR21 U3273 ( .A(a[20]), .B(n2919), .Q(n3546) );
  OAI221 U3274 ( .A(n2924), .B(n2876), .C(n2924), .D(n3548), .Q(n1445) );
  NAND22 U3275 ( .A(n3549), .B(n2850), .Q(n3548) );
  NAND22 U3276 ( .A(n2953), .B(n3550), .Q(n3016) );
  XNR21 U3277 ( .A(a[22]), .B(n2924), .Q(n3550) );
  XNR21 U3278 ( .A(a[22]), .B(n2922), .Q(n3549) );
  OAI221 U3279 ( .A(n2927), .B(n2881), .C(n2927), .D(n3551), .Q(n1444) );
  NAND22 U3280 ( .A(n3552), .B(n2850), .Q(n3551) );
  NAND22 U3281 ( .A(n2950), .B(n3553), .Q(n3018) );
  XNR21 U3282 ( .A(a[24]), .B(n2927), .Q(n3553) );
  XNR21 U3283 ( .A(a[24]), .B(n2924), .Q(n3552) );
  OAI221 U3284 ( .A(n2930), .B(n3020), .C(n2930), .D(n3554), .Q(n1443) );
  NAND22 U3285 ( .A(n3555), .B(n2850), .Q(n3554) );
  NAND22 U3286 ( .A(n2947), .B(n3556), .Q(n3020) );
  XNR21 U3287 ( .A(a[26]), .B(n2930), .Q(n3556) );
  XNR21 U3288 ( .A(a[26]), .B(n2927), .Q(n3555) );
  OAI221 U3289 ( .A(n2933), .B(n2851), .C(n2933), .D(n3557), .Q(n1442) );
  NAND22 U3290 ( .A(n3558), .B(n2850), .Q(n3557) );
  NAND22 U3291 ( .A(n2944), .B(n3559), .Q(n2991) );
  XNR21 U3292 ( .A(a[28]), .B(n2933), .Q(n3559) );
  XNR21 U3293 ( .A(a[28]), .B(n2930), .Q(n3558) );
  OAI221 U3294 ( .A(n2936), .B(n3023), .C(n2936), .D(n3560), .Q(n1441) );
  NAND22 U3295 ( .A(n3561), .B(n2850), .Q(n3560) );
  NAND22 U3296 ( .A(n2940), .B(n3562), .Q(n3023) );
  XNR21 U3297 ( .A(a[30]), .B(n2936), .Q(n3562) );
  XNR21 U3298 ( .A(a[30]), .B(n2933), .Q(n3561) );
endmodule


module Multipliers ( iClk, inRst, iXa, iXb, iYa, iYb, iEn, oX, oY, oReady );
  input [31:0] iXa;
  input [31:0] iXb;
  input [31:0] iYa;
  input [31:0] iYb;
  output [63:0] oX;
  output [63:0] oY;
  input iClk, inRst, iEn;
  output oReady;
  wire   R_STATE__1_, R_STATE__0_, R_XA__31_, R_XA__30_, R_XA__29_, R_XA__28_,
         R_XA__27_, R_XA__26_, R_XA__25_, R_XA__24_, R_XA__23_, R_XA__22_,
         R_XA__21_, R_XA__20_, R_XA__19_, R_XA__18_, R_XA__17_, R_XA__16_,
         R_XA__15_, R_XA__14_, R_XA__13_, R_XA__12_, R_XA__11_, R_XA__10_,
         R_XA__9_, R_XA__8_, R_XA__7_, R_XA__6_, R_XA__5_, R_XA__4_, R_XA__3_,
         R_XA__2_, R_XA__1_, R_XA__0_, R_XB__31_, R_XB__30_, R_XB__29_,
         R_XB__28_, R_XB__27_, R_XB__26_, R_XB__25_, R_XB__24_, R_XB__23_,
         R_XB__22_, R_XB__21_, R_XB__20_, R_XB__19_, R_XB__18_, R_XB__17_,
         R_XB__16_, R_XB__15_, R_XB__14_, R_XB__13_, R_XB__12_, R_XB__11_,
         R_XB__10_, R_XB__9_, R_XB__8_, R_XB__7_, R_XB__6_, R_XB__5_, R_XB__4_,
         R_XB__3_, R_XB__2_, R_XB__1_, R_XB__0_, R_YA__31_, R_YA__30_,
         R_YA__29_, R_YA__28_, R_YA__27_, R_YA__26_, R_YA__25_, R_YA__24_,
         R_YA__23_, R_YA__22_, R_YA__21_, R_YA__20_, R_YA__19_, R_YA__18_,
         R_YA__17_, R_YA__16_, R_YA__15_, R_YA__14_, R_YA__13_, R_YA__12_,
         R_YA__11_, R_YA__10_, R_YA__9_, R_YA__8_, R_YA__7_, R_YA__6_,
         R_YA__5_, R_YA__4_, R_YA__3_, R_YA__2_, R_YA__1_, R_YA__0_, R_YB__31_,
         R_YB__30_, R_YB__29_, R_YB__28_, R_YB__27_, R_YB__26_, R_YB__25_,
         R_YB__24_, R_YB__23_, R_YB__22_, R_YB__21_, R_YB__20_, R_YB__19_,
         R_YB__18_, R_YB__17_, R_YB__16_, R_YB__15_, R_YB__14_, R_YB__13_,
         R_YB__12_, R_YB__11_, R_YB__10_, R_YB__9_, R_YB__8_, R_YB__7_,
         R_YB__6_, R_YB__5_, R_YB__4_, R_YB__3_, R_YB__2_, R_YB__1_, R_YB__0_,
         res_63_, res_62_, res_61_, res_60_, res_59_, res_58_, res_57_,
         res_56_, res_55_, res_54_, res_53_, res_52_, res_51_, res_50_,
         res_49_, res_48_, res_47_, res_46_, res_45_, res_44_, res_43_,
         res_42_, res_41_, res_40_, res_39_, res_38_, res_37_, res_36_,
         res_35_, res_34_, res_33_, res_32_, res_31_, res_30_, res_29_,
         res_28_, res_27_, res_26_, res_25_, res_24_, res_23_, res_22_,
         res_21_, res_20_, res_19_, res_18_, res_17_, res_16_, res_15_,
         res_14_, res_13_, res_12_, res_11_, res_10_, res_9_, res_8_, res_7_,
         res_6_, res_5_, res_4_, res_3_, res_2_, res_1_, res_0_, n262, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998;

  DFEC3 R_reg_STATE__0_ ( .D(n997), .E(n995), .C(iClk), .RN(inRst), .Q(
        R_STATE__0_), .QN(n264) );
  DFC3 R_reg_STATE__1_ ( .D(R_STATE__0_), .C(iClk), .RN(inRst), .Q(R_STATE__1_), .QN(n262) );
  DFEC3 R_reg_YA__31_ ( .D(n971), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__31_) );
  DFC3 R_reg_XA__31_ ( .D(n400), .C(iClk), .RN(inRst), .Q(R_XA__31_) );
  DFEC3 R_reg_YA__30_ ( .D(n963), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__30_) );
  DFC3 R_reg_XA__30_ ( .D(n401), .C(iClk), .RN(inRst), .Q(R_XA__30_) );
  DFEC3 R_reg_YA__29_ ( .D(n955), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__29_) );
  DFC3 R_reg_XA__29_ ( .D(n402), .C(iClk), .RN(inRst), .Q(R_XA__29_) );
  DFEC3 R_reg_YA__28_ ( .D(n947), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__28_) );
  DFC3 R_reg_XA__28_ ( .D(n403), .C(iClk), .RN(inRst), .Q(R_XA__28_) );
  DFEC3 R_reg_YA__27_ ( .D(n939), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__27_) );
  DFC3 R_reg_XA__27_ ( .D(n404), .C(iClk), .RN(inRst), .Q(R_XA__27_) );
  DFEC3 R_reg_YA__26_ ( .D(n931), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__26_) );
  DFC3 R_reg_XA__26_ ( .D(n405), .C(iClk), .RN(inRst), .Q(R_XA__26_) );
  DFEC3 R_reg_YA__25_ ( .D(n923), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__25_) );
  DFC3 R_reg_XA__25_ ( .D(n406), .C(iClk), .RN(inRst), .Q(R_XA__25_) );
  DFEC3 R_reg_YA__24_ ( .D(n915), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__24_) );
  DFC3 R_reg_XA__24_ ( .D(n407), .C(iClk), .RN(inRst), .Q(R_XA__24_) );
  DFEC3 R_reg_YA__23_ ( .D(n907), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__23_) );
  DFC3 R_reg_XA__23_ ( .D(n408), .C(iClk), .RN(inRst), .Q(R_XA__23_) );
  DFEC3 R_reg_YA__22_ ( .D(n899), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__22_) );
  DFC3 R_reg_XA__22_ ( .D(n409), .C(iClk), .RN(inRst), .Q(R_XA__22_) );
  DFEC3 R_reg_YA__21_ ( .D(n891), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__21_) );
  DFC3 R_reg_XA__21_ ( .D(n410), .C(iClk), .RN(inRst), .Q(R_XA__21_) );
  DFEC3 R_reg_YA__20_ ( .D(n883), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__20_) );
  DFC3 R_reg_XA__20_ ( .D(n411), .C(iClk), .RN(inRst), .Q(R_XA__20_) );
  DFEC3 R_reg_YA__19_ ( .D(n875), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__19_) );
  DFC3 R_reg_XA__19_ ( .D(n412), .C(iClk), .RN(inRst), .Q(R_XA__19_) );
  DFEC3 R_reg_YA__18_ ( .D(n867), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__18_) );
  DFC3 R_reg_XA__18_ ( .D(n413), .C(iClk), .RN(inRst), .Q(R_XA__18_) );
  DFEC3 R_reg_YA__17_ ( .D(n859), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__17_) );
  DFC3 R_reg_XA__17_ ( .D(n414), .C(iClk), .RN(inRst), .Q(R_XA__17_) );
  DFEC3 R_reg_YA__16_ ( .D(n851), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__16_) );
  DFC3 R_reg_XA__16_ ( .D(n415), .C(iClk), .RN(inRst), .Q(R_XA__16_) );
  DFEC3 R_reg_YA__15_ ( .D(n843), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__15_) );
  DFC3 R_reg_XA__15_ ( .D(n416), .C(iClk), .RN(inRst), .Q(R_XA__15_) );
  DFEC3 R_reg_YA__14_ ( .D(n835), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__14_) );
  DFC3 R_reg_XA__14_ ( .D(n417), .C(iClk), .RN(inRst), .Q(R_XA__14_) );
  DFEC3 R_reg_YA__13_ ( .D(n827), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__13_) );
  DFC3 R_reg_XA__13_ ( .D(n418), .C(iClk), .RN(inRst), .Q(R_XA__13_) );
  DFEC3 R_reg_YA__12_ ( .D(n819), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__12_) );
  DFC3 R_reg_XA__12_ ( .D(n419), .C(iClk), .RN(inRst), .Q(R_XA__12_) );
  DFEC3 R_reg_YA__11_ ( .D(n811), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__11_) );
  DFC3 R_reg_XA__11_ ( .D(n420), .C(iClk), .RN(inRst), .Q(R_XA__11_) );
  DFEC3 R_reg_YA__10_ ( .D(n803), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__10_) );
  DFC3 R_reg_XA__10_ ( .D(n421), .C(iClk), .RN(inRst), .Q(R_XA__10_) );
  DFEC3 R_reg_YA__9_ ( .D(n795), .E(n985), .C(iClk), .RN(inRst), .Q(R_YA__9_)
         );
  DFC3 R_reg_XA__9_ ( .D(n422), .C(iClk), .RN(inRst), .Q(R_XA__9_) );
  DFEC3 R_reg_YA__8_ ( .D(n787), .E(n986), .C(iClk), .RN(inRst), .Q(R_YA__8_)
         );
  DFC3 R_reg_XA__8_ ( .D(n423), .C(iClk), .RN(inRst), .Q(R_XA__8_) );
  DFEC3 R_reg_YA__7_ ( .D(n779), .E(n987), .C(iClk), .RN(inRst), .Q(R_YA__7_)
         );
  DFC3 R_reg_XA__7_ ( .D(n424), .C(iClk), .RN(inRst), .Q(R_XA__7_) );
  DFEC3 R_reg_YA__6_ ( .D(n771), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__6_)
         );
  DFC3 R_reg_XA__6_ ( .D(n425), .C(iClk), .RN(inRst), .Q(R_XA__6_) );
  DFEC3 R_reg_YA__5_ ( .D(n763), .E(n984), .C(iClk), .RN(inRst), .Q(R_YA__5_)
         );
  DFC3 R_reg_XA__5_ ( .D(n426), .C(iClk), .RN(inRst), .Q(R_XA__5_) );
  DFEC3 R_reg_YA__4_ ( .D(n755), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__4_)
         );
  DFC3 R_reg_XA__4_ ( .D(n427), .C(iClk), .RN(inRst), .Q(R_XA__4_) );
  DFEC3 R_reg_YA__3_ ( .D(n747), .E(n398), .C(iClk), .RN(inRst), .Q(R_YA__3_)
         );
  DFC3 R_reg_XA__3_ ( .D(n428), .C(iClk), .RN(inRst), .Q(R_XA__3_) );
  DFEC3 R_reg_YA__2_ ( .D(n739), .E(n986), .C(iClk), .RN(inRst), .Q(R_YA__2_)
         );
  DFC3 R_reg_XA__2_ ( .D(n429), .C(iClk), .RN(inRst), .Q(R_XA__2_) );
  DFEC3 R_reg_YA__1_ ( .D(n731), .E(n986), .C(iClk), .RN(inRst), .Q(R_YA__1_)
         );
  DFC3 R_reg_XA__1_ ( .D(n430), .C(iClk), .RN(inRst), .Q(R_XA__1_) );
  DFEC3 R_reg_YA__0_ ( .D(n723), .E(n986), .C(iClk), .RN(inRst), .Q(R_YA__0_)
         );
  DFC3 R_reg_XA__0_ ( .D(n431), .C(iClk), .RN(inRst), .Q(R_XA__0_) );
  DFEC3 R_reg_YB__31_ ( .D(n715), .E(n986), .C(iClk), .RN(inRst), .Q(R_YB__31_) );
  DFC3 R_reg_XB__31_ ( .D(n432), .C(iClk), .RN(inRst), .Q(R_XB__31_) );
  DFEC3 R_reg_YB__30_ ( .D(n707), .E(n986), .C(iClk), .RN(inRst), .Q(R_YB__30_) );
  DFC3 R_reg_XB__30_ ( .D(n433), .C(iClk), .RN(inRst), .Q(R_XB__30_) );
  DFEC3 R_reg_YB__29_ ( .D(n699), .E(n986), .C(iClk), .RN(inRst), .Q(R_YB__29_) );
  DFC3 R_reg_XB__29_ ( .D(n434), .C(iClk), .RN(inRst), .Q(R_XB__29_) );
  DFEC3 R_reg_YB__28_ ( .D(n691), .E(n986), .C(iClk), .RN(inRst), .Q(R_YB__28_) );
  DFC3 R_reg_XB__28_ ( .D(n435), .C(iClk), .RN(inRst), .Q(R_XB__28_) );
  DFEC3 R_reg_YB__27_ ( .D(n683), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__27_) );
  DFC3 R_reg_XB__27_ ( .D(n436), .C(iClk), .RN(inRst), .Q(R_XB__27_) );
  DFEC3 R_reg_YB__26_ ( .D(n675), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__26_) );
  DFC3 R_reg_XB__26_ ( .D(n437), .C(iClk), .RN(inRst), .Q(R_XB__26_) );
  DFEC3 R_reg_YB__25_ ( .D(n667), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__25_) );
  DFC3 R_reg_XB__25_ ( .D(n438), .C(iClk), .RN(inRst), .Q(R_XB__25_) );
  DFEC3 R_reg_YB__24_ ( .D(n659), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__24_) );
  DFC3 R_reg_XB__24_ ( .D(n439), .C(iClk), .RN(inRst), .Q(R_XB__24_) );
  DFEC3 R_reg_YB__23_ ( .D(n651), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__23_) );
  DFC3 R_reg_XB__23_ ( .D(n440), .C(iClk), .RN(inRst), .Q(R_XB__23_) );
  DFEC3 R_reg_YB__22_ ( .D(n643), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__22_) );
  DFC3 R_reg_XB__22_ ( .D(n441), .C(iClk), .RN(inRst), .Q(R_XB__22_) );
  DFEC3 R_reg_YB__21_ ( .D(n635), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__21_) );
  DFC3 R_reg_XB__21_ ( .D(n442), .C(iClk), .RN(inRst), .Q(R_XB__21_) );
  DFEC3 R_reg_YB__20_ ( .D(n627), .E(n986), .C(iClk), .RN(inRst), .Q(R_YB__20_) );
  DFC3 R_reg_XB__20_ ( .D(n443), .C(iClk), .RN(inRst), .Q(R_XB__20_) );
  DFEC3 R_reg_YB__19_ ( .D(n619), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__19_) );
  DFC3 R_reg_XB__19_ ( .D(n444), .C(iClk), .RN(inRst), .Q(R_XB__19_) );
  DFEC3 R_reg_YB__18_ ( .D(n611), .E(n984), .C(iClk), .RN(inRst), .Q(R_YB__18_) );
  DFC3 R_reg_XB__18_ ( .D(n445), .C(iClk), .RN(inRst), .Q(R_XB__18_) );
  DFEC3 R_reg_YB__17_ ( .D(n603), .E(n987), .C(iClk), .RN(inRst), .Q(R_YB__17_) );
  DFC3 R_reg_XB__17_ ( .D(n446), .C(iClk), .RN(inRst), .Q(R_XB__17_) );
  DFEC3 R_reg_YB__16_ ( .D(n595), .E(n984), .C(iClk), .RN(inRst), .Q(R_YB__16_) );
  DFC3 R_reg_XB__16_ ( .D(n447), .C(iClk), .RN(inRst), .Q(R_XB__16_) );
  DFEC3 R_reg_YB__15_ ( .D(n587), .E(n984), .C(iClk), .RN(inRst), .Q(R_YB__15_) );
  DFC3 R_reg_XB__15_ ( .D(n448), .C(iClk), .RN(inRst), .Q(R_XB__15_) );
  DFEC3 R_reg_YB__14_ ( .D(n579), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__14_) );
  DFC3 R_reg_XB__14_ ( .D(n449), .C(iClk), .RN(inRst), .Q(R_XB__14_) );
  DFEC3 R_reg_YB__13_ ( .D(n571), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__13_) );
  DFC3 R_reg_XB__13_ ( .D(n450), .C(iClk), .RN(inRst), .Q(R_XB__13_) );
  DFEC3 R_reg_YB__12_ ( .D(n563), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__12_) );
  DFC3 R_reg_XB__12_ ( .D(n451), .C(iClk), .RN(inRst), .Q(R_XB__12_) );
  DFEC3 R_reg_YB__11_ ( .D(n555), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__11_) );
  DFC3 R_reg_XB__11_ ( .D(n452), .C(iClk), .RN(inRst), .Q(R_XB__11_) );
  DFEC3 R_reg_YB__10_ ( .D(n547), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__10_) );
  DFC3 R_reg_XB__10_ ( .D(n453), .C(iClk), .RN(inRst), .Q(R_XB__10_) );
  DFEC3 R_reg_YB__9_ ( .D(n539), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__9_)
         );
  DFC3 R_reg_XB__9_ ( .D(n454), .C(iClk), .RN(inRst), .Q(R_XB__9_) );
  DFEC3 R_reg_YB__8_ ( .D(n531), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__8_)
         );
  DFC3 R_reg_XB__8_ ( .D(n455), .C(iClk), .RN(inRst), .Q(R_XB__8_) );
  DFEC3 R_reg_YB__7_ ( .D(n523), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__7_)
         );
  DFC3 R_reg_XB__7_ ( .D(n456), .C(iClk), .RN(inRst), .Q(R_XB__7_) );
  DFEC3 R_reg_YB__6_ ( .D(n515), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__6_)
         );
  DFC3 R_reg_XB__6_ ( .D(n457), .C(iClk), .RN(inRst), .Q(R_XB__6_) );
  DFEC3 R_reg_YB__5_ ( .D(n507), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__5_)
         );
  DFC3 R_reg_XB__5_ ( .D(n458), .C(iClk), .RN(inRst), .Q(R_XB__5_) );
  DFEC3 R_reg_YB__4_ ( .D(n499), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__4_)
         );
  DFC3 R_reg_XB__4_ ( .D(n459), .C(iClk), .RN(inRst), .Q(R_XB__4_) );
  DFEC3 R_reg_YB__3_ ( .D(n491), .E(n398), .C(iClk), .RN(inRst), .Q(R_YB__3_)
         );
  DFC3 R_reg_XB__3_ ( .D(n460), .C(iClk), .RN(inRst), .Q(R_XB__3_) );
  DFEC3 R_reg_YB__2_ ( .D(n483), .E(n986), .C(iClk), .RN(inRst), .Q(R_YB__2_)
         );
  DFC3 R_reg_XB__2_ ( .D(n461), .C(iClk), .RN(inRst), .Q(R_XB__2_) );
  DFEC3 R_reg_YB__1_ ( .D(n475), .E(n985), .C(iClk), .RN(inRst), .Q(R_YB__1_)
         );
  DFC3 R_reg_XB__1_ ( .D(n462), .C(iClk), .RN(inRst), .Q(R_XB__1_) );
  DFEC3 R_reg_YB__0_ ( .D(n467), .E(n987), .C(iClk), .RN(inRst), .Q(R_YB__0_)
         );
  DFC3 R_reg_XB__0_ ( .D(n463), .C(iClk), .RN(inRst), .Q(R_XB__0_) );
  DFEC3 R_reg_X__63_ ( .D(res_63_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[63])
         );
  DFEC3 R_reg_X__62_ ( .D(res_62_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[62])
         );
  DFEC3 R_reg_X__61_ ( .D(res_61_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[61])
         );
  DFEC3 R_reg_X__60_ ( .D(res_60_), .E(n998), .C(iClk), .RN(inRst), .Q(oX[60])
         );
  DFEC3 R_reg_X__59_ ( .D(res_59_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[59])
         );
  DFEC3 R_reg_X__58_ ( .D(res_58_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[58])
         );
  DFEC3 R_reg_X__57_ ( .D(res_57_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[57])
         );
  DFEC3 R_reg_X__56_ ( .D(res_56_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[56])
         );
  DFEC3 R_reg_X__55_ ( .D(res_55_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[55])
         );
  DFEC3 R_reg_X__54_ ( .D(res_54_), .E(n998), .C(iClk), .RN(inRst), .Q(oX[54])
         );
  DFEC3 R_reg_X__53_ ( .D(res_53_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[53])
         );
  DFEC3 R_reg_X__52_ ( .D(res_52_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[52])
         );
  DFEC3 R_reg_X__51_ ( .D(res_51_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[51])
         );
  DFEC3 R_reg_X__50_ ( .D(res_50_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[50])
         );
  DFEC3 R_reg_X__49_ ( .D(res_49_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[49])
         );
  DFEC3 R_reg_X__48_ ( .D(res_48_), .E(n998), .C(iClk), .RN(inRst), .Q(oX[48])
         );
  DFEC3 R_reg_X__47_ ( .D(res_47_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[47])
         );
  DFEC3 R_reg_X__46_ ( .D(res_46_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[46])
         );
  DFEC3 R_reg_X__45_ ( .D(res_45_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[45])
         );
  DFEC3 R_reg_X__44_ ( .D(res_44_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[44])
         );
  DFEC3 R_reg_X__43_ ( .D(res_43_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[43])
         );
  DFEC3 R_reg_X__42_ ( .D(res_42_), .E(n998), .C(iClk), .RN(inRst), .Q(oX[42])
         );
  DFEC3 R_reg_X__41_ ( .D(res_41_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[41])
         );
  DFEC3 R_reg_X__40_ ( .D(res_40_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[40])
         );
  DFEC3 R_reg_X__39_ ( .D(res_39_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[39])
         );
  DFEC3 R_reg_X__38_ ( .D(res_38_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[38])
         );
  DFEC3 R_reg_X__37_ ( .D(res_37_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[37])
         );
  DFEC3 R_reg_X__36_ ( .D(res_36_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[36])
         );
  DFEC3 R_reg_X__35_ ( .D(res_35_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[35])
         );
  DFEC3 R_reg_X__34_ ( .D(res_34_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[34])
         );
  DFEC3 R_reg_X__33_ ( .D(res_33_), .E(n998), .C(iClk), .RN(inRst), .Q(oX[33])
         );
  DFEC3 R_reg_X__32_ ( .D(res_32_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[32])
         );
  DFEC3 R_reg_X__31_ ( .D(res_31_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[31])
         );
  DFEC3 R_reg_X__30_ ( .D(res_30_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[30])
         );
  DFEC3 R_reg_X__29_ ( .D(res_29_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[29])
         );
  DFEC3 R_reg_X__28_ ( .D(res_28_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[28])
         );
  DFEC3 R_reg_X__27_ ( .D(res_27_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[27])
         );
  DFEC3 R_reg_X__26_ ( .D(res_26_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[26])
         );
  DFEC3 R_reg_X__25_ ( .D(res_25_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[25])
         );
  DFEC3 R_reg_X__24_ ( .D(res_24_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[24])
         );
  DFEC3 R_reg_X__23_ ( .D(res_23_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[23])
         );
  DFEC3 R_reg_X__22_ ( .D(res_22_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[22])
         );
  DFEC3 R_reg_X__21_ ( .D(res_21_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[21])
         );
  DFEC3 R_reg_X__20_ ( .D(res_20_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[20])
         );
  DFEC3 R_reg_X__19_ ( .D(res_19_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[19])
         );
  DFEC3 R_reg_X__18_ ( .D(res_18_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[18])
         );
  DFEC3 R_reg_X__17_ ( .D(res_17_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[17])
         );
  DFEC3 R_reg_X__16_ ( .D(res_16_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[16])
         );
  DFEC3 R_reg_X__15_ ( .D(res_15_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[15])
         );
  DFEC3 R_reg_X__14_ ( .D(res_14_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[14])
         );
  DFEC3 R_reg_X__13_ ( .D(res_13_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[13])
         );
  DFEC3 R_reg_X__12_ ( .D(res_12_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[12])
         );
  DFEC3 R_reg_X__11_ ( .D(res_11_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[11])
         );
  DFEC3 R_reg_X__10_ ( .D(res_10_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[10])
         );
  DFEC3 R_reg_X__9_ ( .D(res_9_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[9]) );
  DFEC3 R_reg_X__8_ ( .D(res_8_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[8]) );
  DFEC3 R_reg_X__7_ ( .D(res_7_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[7]) );
  DFEC3 R_reg_X__6_ ( .D(res_6_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[6]) );
  DFEC3 R_reg_X__5_ ( .D(res_5_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[5]) );
  DFEC3 R_reg_X__4_ ( .D(res_4_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[4]) );
  DFEC3 R_reg_X__3_ ( .D(res_3_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[3]) );
  DFEC3 R_reg_X__2_ ( .D(res_2_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[2]) );
  DFEC3 R_reg_X__1_ ( .D(res_1_), .E(n982), .C(iClk), .RN(inRst), .Q(oX[1]) );
  DFEC3 R_reg_X__0_ ( .D(res_0_), .E(n983), .C(iClk), .RN(inRst), .Q(oX[0]) );
  DFEC3 R_reg_Y__63_ ( .D(res_63_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[63])
         );
  DFEC3 R_reg_Y__62_ ( .D(res_62_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[62])
         );
  DFEC3 R_reg_Y__61_ ( .D(res_61_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[61])
         );
  DFEC3 R_reg_Y__60_ ( .D(res_60_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[60])
         );
  DFEC3 R_reg_Y__59_ ( .D(res_59_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[59])
         );
  DFEC3 R_reg_Y__58_ ( .D(res_58_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[58])
         );
  DFEC3 R_reg_Y__57_ ( .D(res_57_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[57])
         );
  DFEC3 R_reg_Y__56_ ( .D(res_56_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[56])
         );
  DFEC3 R_reg_Y__55_ ( .D(res_55_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[55])
         );
  DFEC3 R_reg_Y__54_ ( .D(res_54_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[54])
         );
  DFEC3 R_reg_Y__53_ ( .D(res_53_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[53])
         );
  DFEC3 R_reg_Y__52_ ( .D(res_52_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[52])
         );
  DFEC3 R_reg_Y__51_ ( .D(res_51_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[51])
         );
  DFEC3 R_reg_Y__50_ ( .D(res_50_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[50])
         );
  DFEC3 R_reg_Y__49_ ( .D(res_49_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[49])
         );
  DFEC3 R_reg_Y__48_ ( .D(res_48_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[48])
         );
  DFEC3 R_reg_Y__47_ ( .D(res_47_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[47])
         );
  DFEC3 R_reg_Y__46_ ( .D(res_46_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[46])
         );
  DFEC3 R_reg_Y__45_ ( .D(res_45_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[45])
         );
  DFEC3 R_reg_Y__44_ ( .D(res_44_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[44])
         );
  DFEC3 R_reg_Y__43_ ( .D(res_43_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[43])
         );
  DFEC3 R_reg_Y__42_ ( .D(res_42_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[42])
         );
  DFEC3 R_reg_Y__41_ ( .D(res_41_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[41])
         );
  DFEC3 R_reg_Y__40_ ( .D(res_40_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[40])
         );
  DFEC3 R_reg_Y__39_ ( .D(res_39_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[39])
         );
  DFEC3 R_reg_Y__38_ ( .D(res_38_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[38])
         );
  DFEC3 R_reg_Y__37_ ( .D(res_37_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[37])
         );
  DFEC3 R_reg_Y__36_ ( .D(res_36_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[36])
         );
  DFEC3 R_reg_Y__35_ ( .D(res_35_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[35])
         );
  DFEC3 R_reg_Y__34_ ( .D(res_34_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[34])
         );
  DFEC3 R_reg_Y__33_ ( .D(res_33_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[33])
         );
  DFEC3 R_reg_Y__32_ ( .D(res_32_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[32])
         );
  DFEC3 R_reg_Y__31_ ( .D(res_31_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[31])
         );
  DFEC3 R_reg_Y__30_ ( .D(res_30_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[30])
         );
  DFEC3 R_reg_Y__29_ ( .D(res_29_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[29])
         );
  DFEC3 R_reg_Y__28_ ( .D(res_28_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[28])
         );
  DFEC3 R_reg_Y__27_ ( .D(res_27_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[27])
         );
  DFEC3 R_reg_Y__26_ ( .D(res_26_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[26])
         );
  DFEC3 R_reg_Y__25_ ( .D(res_25_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[25])
         );
  DFEC3 R_reg_Y__24_ ( .D(res_24_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[24])
         );
  DFEC3 R_reg_Y__23_ ( .D(res_23_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[23])
         );
  DFEC3 R_reg_Y__22_ ( .D(res_22_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[22])
         );
  DFEC3 R_reg_Y__21_ ( .D(res_21_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[21])
         );
  DFEC3 R_reg_Y__20_ ( .D(res_20_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[20])
         );
  DFEC3 R_reg_Y__19_ ( .D(res_19_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[19])
         );
  DFEC3 R_reg_Y__18_ ( .D(res_18_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[18])
         );
  DFEC3 R_reg_Y__17_ ( .D(res_17_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[17])
         );
  DFEC3 R_reg_Y__16_ ( .D(res_16_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[16])
         );
  DFEC3 R_reg_Y__15_ ( .D(res_15_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[15])
         );
  DFEC3 R_reg_Y__14_ ( .D(res_14_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[14])
         );
  DFEC3 R_reg_Y__13_ ( .D(res_13_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[13])
         );
  DFEC3 R_reg_Y__12_ ( .D(res_12_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[12])
         );
  DFEC3 R_reg_Y__11_ ( .D(res_11_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[11])
         );
  DFEC3 R_reg_Y__10_ ( .D(res_10_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[10])
         );
  DFEC3 R_reg_Y__9_ ( .D(res_9_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[9]) );
  DFEC3 R_reg_Y__8_ ( .D(res_8_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[8]) );
  DFEC3 R_reg_Y__7_ ( .D(res_7_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[7]) );
  DFEC3 R_reg_Y__6_ ( .D(res_6_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[6]) );
  DFEC3 R_reg_Y__5_ ( .D(res_5_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[5]) );
  DFEC3 R_reg_Y__4_ ( .D(res_4_), .E(n979), .C(iClk), .RN(inRst), .Q(oY[4]) );
  DFEC3 R_reg_Y__3_ ( .D(res_3_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[3]) );
  DFEC3 R_reg_Y__2_ ( .D(res_2_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[2]) );
  DFEC3 R_reg_Y__1_ ( .D(res_1_), .E(n981), .C(iClk), .RN(inRst), .Q(oY[1]) );
  DFEC3 R_reg_Y__0_ ( .D(res_0_), .E(n980), .C(iClk), .RN(inRst), .Q(oY[0]) );
  DFC3 R_reg_READY_ ( .D(n979), .C(iClk), .RN(inRst), .Q(oReady) );
  Multipliers_DW_mult_tc_0 mult_68 ( .a({R_XA__31_, R_XA__30_, R_XA__29_, 
        R_XA__28_, R_XA__27_, R_XA__26_, R_XA__25_, R_XA__24_, R_XA__23_, 
        R_XA__22_, R_XA__21_, R_XA__20_, R_XA__19_, R_XA__18_, R_XA__17_, 
        R_XA__16_, R_XA__15_, R_XA__14_, R_XA__13_, R_XA__12_, R_XA__11_, 
        R_XA__10_, R_XA__9_, R_XA__8_, R_XA__7_, R_XA__6_, R_XA__5_, R_XA__4_, 
        R_XA__3_, R_XA__2_, R_XA__1_, R_XA__0_}), .b({R_XB__31_, R_XB__30_, 
        R_XB__29_, R_XB__28_, R_XB__27_, R_XB__26_, R_XB__25_, R_XB__24_, 
        R_XB__23_, R_XB__22_, R_XB__21_, R_XB__20_, R_XB__19_, R_XB__18_, 
        R_XB__17_, R_XB__16_, R_XB__15_, R_XB__14_, R_XB__13_, R_XB__12_, 
        R_XB__11_, R_XB__10_, R_XB__9_, R_XB__8_, R_XB__7_, R_XB__6_, R_XB__5_, 
        R_XB__4_, R_XB__3_, R_XB__2_, R_XB__1_, R_XB__0_}), .product({res_63_, 
        res_62_, res_61_, res_60_, res_59_, res_58_, res_57_, res_56_, res_55_, 
        res_54_, res_53_, res_52_, res_51_, res_50_, res_49_, res_48_, res_47_, 
        res_46_, res_45_, res_44_, res_43_, res_42_, res_41_, res_40_, res_39_, 
        res_38_, res_37_, res_36_, res_35_, res_34_, res_33_, res_32_, res_31_, 
        res_30_, res_29_, res_28_, res_27_, res_26_, res_25_, res_24_, res_23_, 
        res_22_, res_21_, res_20_, res_19_, res_18_, res_17_, res_16_, res_15_, 
        res_14_, res_13_, res_12_, res_11_, res_10_, res_9_, res_8_, res_7_, 
        res_6_, res_5_, res_4_, res_3_, res_2_, res_1_, res_0_}) );
  NOR22 U207 ( .A(n262), .B(R_STATE__0_), .Q(n996) );
  NOR22 U208 ( .A(n998), .B(n269), .Q(n398) );
  NOR22 U209 ( .A(n262), .B(R_STATE__0_), .Q(n981) );
  NOR22 U210 ( .A(R_STATE__0_), .B(R_STATE__1_), .Q(n997) );
  CLKBU6 U211 ( .A(n465), .Q(n464) );
  CLKBU6 U212 ( .A(n466), .Q(n465) );
  CLKBU6 U213 ( .A(iXb[0]), .Q(n466) );
  CLKBU6 U214 ( .A(n468), .Q(n467) );
  CLKBU6 U215 ( .A(n469), .Q(n468) );
  CLKBU6 U216 ( .A(n470), .Q(n469) );
  CLKBU6 U217 ( .A(n471), .Q(n470) );
  CLKBU6 U218 ( .A(iYb[0]), .Q(n471) );
  CLKBU6 U219 ( .A(n473), .Q(n472) );
  CLKBU6 U220 ( .A(n474), .Q(n473) );
  CLKBU6 U221 ( .A(iXb[1]), .Q(n474) );
  CLKBU6 U222 ( .A(n476), .Q(n475) );
  CLKBU6 U223 ( .A(n477), .Q(n476) );
  CLKBU6 U224 ( .A(n478), .Q(n477) );
  CLKBU6 U225 ( .A(n479), .Q(n478) );
  CLKBU6 U226 ( .A(iYb[1]), .Q(n479) );
  CLKBU6 U227 ( .A(n481), .Q(n480) );
  CLKBU6 U228 ( .A(n482), .Q(n481) );
  CLKBU6 U229 ( .A(iXb[2]), .Q(n482) );
  CLKBU6 U230 ( .A(n484), .Q(n483) );
  CLKBU6 U231 ( .A(n485), .Q(n484) );
  CLKBU6 U232 ( .A(n486), .Q(n485) );
  CLKBU6 U233 ( .A(n487), .Q(n486) );
  CLKBU6 U234 ( .A(iYb[2]), .Q(n487) );
  CLKBU6 U235 ( .A(n489), .Q(n488) );
  CLKBU6 U236 ( .A(n490), .Q(n489) );
  CLKBU6 U237 ( .A(iXb[3]), .Q(n490) );
  CLKBU6 U238 ( .A(n492), .Q(n491) );
  CLKBU6 U239 ( .A(n493), .Q(n492) );
  CLKBU6 U240 ( .A(n494), .Q(n493) );
  CLKBU6 U241 ( .A(n495), .Q(n494) );
  CLKBU6 U242 ( .A(iYb[3]), .Q(n495) );
  CLKBU6 U243 ( .A(n497), .Q(n496) );
  CLKBU6 U244 ( .A(n498), .Q(n497) );
  CLKBU6 U245 ( .A(iXb[4]), .Q(n498) );
  CLKBU6 U246 ( .A(n500), .Q(n499) );
  CLKBU6 U247 ( .A(n501), .Q(n500) );
  CLKBU6 U248 ( .A(n502), .Q(n501) );
  CLKBU6 U249 ( .A(n503), .Q(n502) );
  CLKBU6 U250 ( .A(iYb[4]), .Q(n503) );
  CLKBU6 U251 ( .A(n505), .Q(n504) );
  CLKBU6 U252 ( .A(n506), .Q(n505) );
  CLKBU6 U253 ( .A(iXb[5]), .Q(n506) );
  CLKBU6 U254 ( .A(n508), .Q(n507) );
  CLKBU6 U255 ( .A(n509), .Q(n508) );
  CLKBU6 U256 ( .A(n510), .Q(n509) );
  CLKBU6 U257 ( .A(n511), .Q(n510) );
  CLKBU6 U258 ( .A(iYb[5]), .Q(n511) );
  CLKBU6 U259 ( .A(n513), .Q(n512) );
  CLKBU6 U260 ( .A(n514), .Q(n513) );
  CLKBU6 U261 ( .A(iXb[6]), .Q(n514) );
  CLKBU6 U262 ( .A(n516), .Q(n515) );
  CLKBU6 U263 ( .A(n517), .Q(n516) );
  CLKBU6 U264 ( .A(n518), .Q(n517) );
  CLKBU6 U265 ( .A(n519), .Q(n518) );
  CLKBU6 U266 ( .A(iYb[6]), .Q(n519) );
  CLKBU6 U267 ( .A(n521), .Q(n520) );
  CLKBU6 U268 ( .A(n522), .Q(n521) );
  CLKBU6 U269 ( .A(iXb[7]), .Q(n522) );
  CLKBU6 U270 ( .A(n524), .Q(n523) );
  CLKBU6 U271 ( .A(n525), .Q(n524) );
  CLKBU6 U272 ( .A(n526), .Q(n525) );
  CLKBU6 U273 ( .A(n527), .Q(n526) );
  CLKBU6 U274 ( .A(iYb[7]), .Q(n527) );
  CLKBU6 U275 ( .A(n529), .Q(n528) );
  CLKBU6 U276 ( .A(n530), .Q(n529) );
  CLKBU6 U277 ( .A(iXb[8]), .Q(n530) );
  CLKBU6 U278 ( .A(n532), .Q(n531) );
  CLKBU6 U279 ( .A(n533), .Q(n532) );
  CLKBU6 U280 ( .A(n534), .Q(n533) );
  CLKBU6 U281 ( .A(n535), .Q(n534) );
  CLKBU6 U282 ( .A(iYb[8]), .Q(n535) );
  CLKBU6 U283 ( .A(n537), .Q(n536) );
  CLKBU6 U284 ( .A(n538), .Q(n537) );
  CLKBU6 U285 ( .A(iXb[9]), .Q(n538) );
  CLKBU6 U286 ( .A(n540), .Q(n539) );
  CLKBU6 U287 ( .A(n541), .Q(n540) );
  CLKBU6 U288 ( .A(n542), .Q(n541) );
  CLKBU6 U289 ( .A(n543), .Q(n542) );
  CLKBU6 U290 ( .A(iYb[9]), .Q(n543) );
  CLKBU6 U291 ( .A(n545), .Q(n544) );
  CLKBU6 U292 ( .A(n546), .Q(n545) );
  CLKBU6 U293 ( .A(iXb[10]), .Q(n546) );
  CLKBU6 U294 ( .A(n548), .Q(n547) );
  CLKBU6 U295 ( .A(n549), .Q(n548) );
  CLKBU6 U296 ( .A(n550), .Q(n549) );
  CLKBU6 U297 ( .A(n551), .Q(n550) );
  CLKBU6 U298 ( .A(iYb[10]), .Q(n551) );
  CLKBU6 U299 ( .A(n553), .Q(n552) );
  CLKBU6 U300 ( .A(n554), .Q(n553) );
  CLKBU6 U301 ( .A(iXb[11]), .Q(n554) );
  CLKBU6 U302 ( .A(n556), .Q(n555) );
  CLKBU6 U303 ( .A(n557), .Q(n556) );
  CLKBU6 U304 ( .A(n558), .Q(n557) );
  CLKBU6 U305 ( .A(n559), .Q(n558) );
  CLKBU6 U306 ( .A(iYb[11]), .Q(n559) );
  CLKBU6 U307 ( .A(n561), .Q(n560) );
  CLKBU6 U308 ( .A(n562), .Q(n561) );
  CLKBU6 U309 ( .A(iXb[12]), .Q(n562) );
  CLKBU6 U310 ( .A(n564), .Q(n563) );
  CLKBU6 U311 ( .A(n565), .Q(n564) );
  CLKBU6 U312 ( .A(n566), .Q(n565) );
  CLKBU6 U313 ( .A(n567), .Q(n566) );
  CLKBU6 U314 ( .A(iYb[12]), .Q(n567) );
  CLKBU6 U315 ( .A(n569), .Q(n568) );
  CLKBU6 U316 ( .A(n570), .Q(n569) );
  CLKBU6 U317 ( .A(iXb[13]), .Q(n570) );
  CLKBU6 U318 ( .A(n572), .Q(n571) );
  CLKBU6 U319 ( .A(n573), .Q(n572) );
  CLKBU6 U320 ( .A(n574), .Q(n573) );
  CLKBU6 U321 ( .A(n575), .Q(n574) );
  CLKBU6 U322 ( .A(iYb[13]), .Q(n575) );
  CLKBU6 U323 ( .A(n577), .Q(n576) );
  CLKBU6 U324 ( .A(n578), .Q(n577) );
  CLKBU6 U325 ( .A(iXb[14]), .Q(n578) );
  CLKBU6 U326 ( .A(n580), .Q(n579) );
  CLKBU6 U327 ( .A(n581), .Q(n580) );
  CLKBU6 U328 ( .A(n582), .Q(n581) );
  CLKBU6 U329 ( .A(n583), .Q(n582) );
  CLKBU6 U330 ( .A(iYb[14]), .Q(n583) );
  CLKBU6 U331 ( .A(n585), .Q(n584) );
  CLKBU6 U332 ( .A(n586), .Q(n585) );
  CLKBU6 U333 ( .A(iXb[15]), .Q(n586) );
  CLKBU6 U334 ( .A(n588), .Q(n587) );
  CLKBU6 U335 ( .A(n589), .Q(n588) );
  CLKBU6 U336 ( .A(n590), .Q(n589) );
  CLKBU6 U337 ( .A(n591), .Q(n590) );
  CLKBU6 U338 ( .A(iYb[15]), .Q(n591) );
  CLKBU6 U339 ( .A(n593), .Q(n592) );
  CLKBU6 U340 ( .A(n594), .Q(n593) );
  CLKBU6 U341 ( .A(iXb[16]), .Q(n594) );
  CLKBU6 U342 ( .A(n596), .Q(n595) );
  CLKBU6 U343 ( .A(n597), .Q(n596) );
  CLKBU6 U344 ( .A(n598), .Q(n597) );
  CLKBU6 U345 ( .A(n599), .Q(n598) );
  CLKBU6 U346 ( .A(iYb[16]), .Q(n599) );
  CLKBU6 U347 ( .A(n601), .Q(n600) );
  CLKBU6 U348 ( .A(n602), .Q(n601) );
  CLKBU6 U349 ( .A(iXb[17]), .Q(n602) );
  CLKBU6 U350 ( .A(n604), .Q(n603) );
  CLKBU6 U351 ( .A(n605), .Q(n604) );
  CLKBU6 U352 ( .A(n606), .Q(n605) );
  CLKBU6 U353 ( .A(n607), .Q(n606) );
  CLKBU6 U354 ( .A(iYb[17]), .Q(n607) );
  CLKBU6 U355 ( .A(n609), .Q(n608) );
  CLKBU6 U356 ( .A(n610), .Q(n609) );
  CLKBU6 U357 ( .A(iXb[18]), .Q(n610) );
  CLKBU6 U358 ( .A(n612), .Q(n611) );
  CLKBU6 U359 ( .A(n613), .Q(n612) );
  CLKBU6 U360 ( .A(n614), .Q(n613) );
  CLKBU6 U361 ( .A(n615), .Q(n614) );
  CLKBU6 U362 ( .A(iYb[18]), .Q(n615) );
  CLKBU6 U363 ( .A(n617), .Q(n616) );
  CLKBU6 U364 ( .A(n618), .Q(n617) );
  CLKBU6 U365 ( .A(iXb[19]), .Q(n618) );
  CLKBU6 U366 ( .A(n620), .Q(n619) );
  CLKBU6 U367 ( .A(n621), .Q(n620) );
  CLKBU6 U368 ( .A(n622), .Q(n621) );
  CLKBU6 U369 ( .A(n623), .Q(n622) );
  CLKBU6 U370 ( .A(iYb[19]), .Q(n623) );
  CLKBU6 U371 ( .A(n625), .Q(n624) );
  CLKBU6 U372 ( .A(n626), .Q(n625) );
  CLKBU6 U373 ( .A(iXb[20]), .Q(n626) );
  CLKBU6 U374 ( .A(n628), .Q(n627) );
  CLKBU6 U375 ( .A(n629), .Q(n628) );
  CLKBU6 U376 ( .A(n630), .Q(n629) );
  CLKBU6 U377 ( .A(n631), .Q(n630) );
  CLKBU6 U378 ( .A(iYb[20]), .Q(n631) );
  CLKBU6 U379 ( .A(n633), .Q(n632) );
  CLKBU6 U380 ( .A(n634), .Q(n633) );
  CLKBU6 U381 ( .A(iXb[21]), .Q(n634) );
  CLKBU6 U382 ( .A(n636), .Q(n635) );
  CLKBU6 U383 ( .A(n637), .Q(n636) );
  CLKBU6 U384 ( .A(n638), .Q(n637) );
  CLKBU6 U385 ( .A(n639), .Q(n638) );
  CLKBU6 U386 ( .A(iYb[21]), .Q(n639) );
  CLKBU6 U387 ( .A(n641), .Q(n640) );
  CLKBU6 U388 ( .A(n642), .Q(n641) );
  CLKBU6 U389 ( .A(iXb[22]), .Q(n642) );
  CLKBU6 U390 ( .A(n644), .Q(n643) );
  CLKBU6 U391 ( .A(n645), .Q(n644) );
  CLKBU6 U392 ( .A(n646), .Q(n645) );
  CLKBU6 U393 ( .A(n647), .Q(n646) );
  CLKBU6 U394 ( .A(iYb[22]), .Q(n647) );
  CLKBU6 U395 ( .A(n649), .Q(n648) );
  CLKBU6 U396 ( .A(n650), .Q(n649) );
  CLKBU6 U397 ( .A(iXb[23]), .Q(n650) );
  CLKBU6 U398 ( .A(n652), .Q(n651) );
  CLKBU6 U399 ( .A(n653), .Q(n652) );
  CLKBU6 U400 ( .A(n654), .Q(n653) );
  CLKBU6 U401 ( .A(n655), .Q(n654) );
  CLKBU6 U402 ( .A(iYb[23]), .Q(n655) );
  CLKBU6 U403 ( .A(n657), .Q(n656) );
  CLKBU6 U404 ( .A(n658), .Q(n657) );
  CLKBU6 U405 ( .A(iXb[24]), .Q(n658) );
  CLKBU6 U406 ( .A(n660), .Q(n659) );
  CLKBU6 U407 ( .A(n661), .Q(n660) );
  CLKBU6 U408 ( .A(n662), .Q(n661) );
  CLKBU6 U409 ( .A(n663), .Q(n662) );
  CLKBU6 U410 ( .A(iYb[24]), .Q(n663) );
  CLKBU6 U411 ( .A(n665), .Q(n664) );
  CLKBU6 U412 ( .A(n666), .Q(n665) );
  CLKBU6 U413 ( .A(iXb[25]), .Q(n666) );
  CLKBU6 U414 ( .A(n668), .Q(n667) );
  CLKBU6 U415 ( .A(n669), .Q(n668) );
  CLKBU6 U416 ( .A(n670), .Q(n669) );
  CLKBU6 U417 ( .A(n671), .Q(n670) );
  CLKBU6 U418 ( .A(iYb[25]), .Q(n671) );
  CLKBU6 U419 ( .A(n673), .Q(n672) );
  CLKBU6 U420 ( .A(n674), .Q(n673) );
  CLKBU6 U421 ( .A(iXb[26]), .Q(n674) );
  CLKBU6 U422 ( .A(n676), .Q(n675) );
  CLKBU6 U423 ( .A(n677), .Q(n676) );
  CLKBU6 U424 ( .A(n678), .Q(n677) );
  CLKBU6 U425 ( .A(n679), .Q(n678) );
  CLKBU6 U426 ( .A(iYb[26]), .Q(n679) );
  CLKBU6 U427 ( .A(n681), .Q(n680) );
  CLKBU6 U428 ( .A(n682), .Q(n681) );
  CLKBU6 U429 ( .A(iXb[27]), .Q(n682) );
  CLKBU6 U430 ( .A(n684), .Q(n683) );
  CLKBU6 U431 ( .A(n685), .Q(n684) );
  CLKBU6 U432 ( .A(n686), .Q(n685) );
  CLKBU6 U433 ( .A(n687), .Q(n686) );
  CLKBU6 U434 ( .A(iYb[27]), .Q(n687) );
  CLKBU6 U435 ( .A(n689), .Q(n688) );
  CLKBU6 U436 ( .A(n690), .Q(n689) );
  CLKBU6 U437 ( .A(iXb[28]), .Q(n690) );
  CLKBU6 U438 ( .A(n692), .Q(n691) );
  CLKBU6 U439 ( .A(n693), .Q(n692) );
  CLKBU6 U440 ( .A(n694), .Q(n693) );
  CLKBU6 U441 ( .A(n695), .Q(n694) );
  CLKBU6 U442 ( .A(iYb[28]), .Q(n695) );
  CLKBU6 U443 ( .A(n697), .Q(n696) );
  CLKBU6 U444 ( .A(n698), .Q(n697) );
  CLKBU6 U445 ( .A(iXb[29]), .Q(n698) );
  CLKBU6 U446 ( .A(n700), .Q(n699) );
  CLKBU6 U447 ( .A(n701), .Q(n700) );
  CLKBU6 U448 ( .A(n702), .Q(n701) );
  CLKBU6 U449 ( .A(n703), .Q(n702) );
  CLKBU6 U450 ( .A(iYb[29]), .Q(n703) );
  CLKBU6 U451 ( .A(n705), .Q(n704) );
  CLKBU6 U452 ( .A(n706), .Q(n705) );
  CLKBU6 U453 ( .A(iXb[30]), .Q(n706) );
  CLKBU6 U454 ( .A(n708), .Q(n707) );
  CLKBU6 U455 ( .A(n709), .Q(n708) );
  CLKBU6 U456 ( .A(n710), .Q(n709) );
  CLKBU6 U457 ( .A(n711), .Q(n710) );
  CLKBU6 U458 ( .A(iYb[30]), .Q(n711) );
  CLKBU6 U459 ( .A(n713), .Q(n712) );
  CLKBU6 U460 ( .A(n714), .Q(n713) );
  CLKBU6 U461 ( .A(iXb[31]), .Q(n714) );
  CLKBU6 U462 ( .A(n716), .Q(n715) );
  CLKBU6 U463 ( .A(n717), .Q(n716) );
  CLKBU6 U464 ( .A(n718), .Q(n717) );
  CLKBU6 U465 ( .A(n719), .Q(n718) );
  CLKBU6 U466 ( .A(iYb[31]), .Q(n719) );
  CLKBU6 U467 ( .A(n721), .Q(n720) );
  CLKBU6 U468 ( .A(n722), .Q(n721) );
  CLKBU6 U469 ( .A(iXa[0]), .Q(n722) );
  CLKBU6 U470 ( .A(n724), .Q(n723) );
  CLKBU6 U471 ( .A(n725), .Q(n724) );
  CLKBU6 U472 ( .A(n726), .Q(n725) );
  CLKBU6 U473 ( .A(n727), .Q(n726) );
  CLKBU6 U474 ( .A(iYa[0]), .Q(n727) );
  CLKBU6 U475 ( .A(n729), .Q(n728) );
  CLKBU6 U476 ( .A(n730), .Q(n729) );
  CLKBU6 U477 ( .A(iXa[1]), .Q(n730) );
  CLKBU6 U478 ( .A(n732), .Q(n731) );
  CLKBU6 U479 ( .A(n733), .Q(n732) );
  CLKBU6 U480 ( .A(n734), .Q(n733) );
  CLKBU6 U481 ( .A(n735), .Q(n734) );
  CLKBU6 U482 ( .A(iYa[1]), .Q(n735) );
  CLKBU6 U483 ( .A(n737), .Q(n736) );
  CLKBU6 U484 ( .A(n738), .Q(n737) );
  CLKBU6 U485 ( .A(iXa[2]), .Q(n738) );
  CLKBU6 U486 ( .A(n740), .Q(n739) );
  CLKBU6 U487 ( .A(n741), .Q(n740) );
  CLKBU6 U488 ( .A(n742), .Q(n741) );
  CLKBU6 U489 ( .A(n743), .Q(n742) );
  CLKBU6 U490 ( .A(iYa[2]), .Q(n743) );
  CLKBU6 U491 ( .A(n745), .Q(n744) );
  CLKBU6 U492 ( .A(n746), .Q(n745) );
  CLKBU6 U493 ( .A(iXa[3]), .Q(n746) );
  CLKBU6 U494 ( .A(n748), .Q(n747) );
  CLKBU6 U495 ( .A(n749), .Q(n748) );
  CLKBU6 U496 ( .A(n750), .Q(n749) );
  CLKBU6 U497 ( .A(n751), .Q(n750) );
  CLKBU6 U498 ( .A(iYa[3]), .Q(n751) );
  CLKBU6 U499 ( .A(n753), .Q(n752) );
  CLKBU6 U500 ( .A(n754), .Q(n753) );
  CLKBU6 U501 ( .A(iXa[4]), .Q(n754) );
  CLKBU6 U502 ( .A(n756), .Q(n755) );
  CLKBU6 U503 ( .A(n757), .Q(n756) );
  CLKBU6 U504 ( .A(n758), .Q(n757) );
  CLKBU6 U505 ( .A(n759), .Q(n758) );
  CLKBU6 U506 ( .A(iYa[4]), .Q(n759) );
  CLKBU6 U507 ( .A(n761), .Q(n760) );
  CLKBU6 U508 ( .A(n762), .Q(n761) );
  CLKBU6 U509 ( .A(iXa[5]), .Q(n762) );
  CLKBU6 U510 ( .A(n764), .Q(n763) );
  CLKBU6 U511 ( .A(n765), .Q(n764) );
  CLKBU6 U512 ( .A(n766), .Q(n765) );
  CLKBU6 U513 ( .A(n767), .Q(n766) );
  CLKBU6 U514 ( .A(iYa[5]), .Q(n767) );
  CLKBU6 U515 ( .A(n769), .Q(n768) );
  CLKBU6 U516 ( .A(n770), .Q(n769) );
  CLKBU6 U517 ( .A(iXa[6]), .Q(n770) );
  CLKBU6 U518 ( .A(n772), .Q(n771) );
  CLKBU6 U519 ( .A(n773), .Q(n772) );
  CLKBU6 U520 ( .A(n774), .Q(n773) );
  CLKBU6 U521 ( .A(n775), .Q(n774) );
  CLKBU6 U522 ( .A(iYa[6]), .Q(n775) );
  CLKBU6 U523 ( .A(n777), .Q(n776) );
  CLKBU6 U524 ( .A(n778), .Q(n777) );
  CLKBU6 U525 ( .A(iXa[7]), .Q(n778) );
  CLKBU6 U526 ( .A(n780), .Q(n779) );
  CLKBU6 U527 ( .A(n781), .Q(n780) );
  CLKBU6 U528 ( .A(n782), .Q(n781) );
  CLKBU6 U529 ( .A(n783), .Q(n782) );
  CLKBU6 U530 ( .A(iYa[7]), .Q(n783) );
  CLKBU6 U531 ( .A(n785), .Q(n784) );
  CLKBU6 U532 ( .A(n786), .Q(n785) );
  CLKBU6 U533 ( .A(iXa[8]), .Q(n786) );
  CLKBU6 U534 ( .A(n788), .Q(n787) );
  CLKBU6 U535 ( .A(n789), .Q(n788) );
  CLKBU6 U536 ( .A(n790), .Q(n789) );
  CLKBU6 U537 ( .A(n791), .Q(n790) );
  CLKBU6 U538 ( .A(iYa[8]), .Q(n791) );
  CLKBU6 U539 ( .A(n793), .Q(n792) );
  CLKBU6 U540 ( .A(n794), .Q(n793) );
  CLKBU6 U541 ( .A(iXa[9]), .Q(n794) );
  CLKBU6 U542 ( .A(n796), .Q(n795) );
  CLKBU6 U543 ( .A(n797), .Q(n796) );
  CLKBU6 U544 ( .A(n798), .Q(n797) );
  CLKBU6 U545 ( .A(n799), .Q(n798) );
  CLKBU6 U546 ( .A(iYa[9]), .Q(n799) );
  CLKBU6 U547 ( .A(n801), .Q(n800) );
  CLKBU6 U548 ( .A(n802), .Q(n801) );
  CLKBU6 U549 ( .A(iXa[10]), .Q(n802) );
  CLKBU6 U550 ( .A(n804), .Q(n803) );
  CLKBU6 U551 ( .A(n805), .Q(n804) );
  CLKBU6 U552 ( .A(n806), .Q(n805) );
  CLKBU6 U553 ( .A(n807), .Q(n806) );
  CLKBU6 U554 ( .A(iYa[10]), .Q(n807) );
  CLKBU6 U555 ( .A(n809), .Q(n808) );
  CLKBU6 U556 ( .A(n810), .Q(n809) );
  CLKBU6 U557 ( .A(iXa[11]), .Q(n810) );
  CLKBU6 U558 ( .A(n812), .Q(n811) );
  CLKBU6 U559 ( .A(n813), .Q(n812) );
  CLKBU6 U560 ( .A(n814), .Q(n813) );
  CLKBU6 U561 ( .A(n815), .Q(n814) );
  CLKBU6 U562 ( .A(iYa[11]), .Q(n815) );
  CLKBU6 U563 ( .A(n817), .Q(n816) );
  CLKBU6 U564 ( .A(n818), .Q(n817) );
  CLKBU6 U565 ( .A(iXa[12]), .Q(n818) );
  CLKBU6 U566 ( .A(n820), .Q(n819) );
  CLKBU6 U567 ( .A(n821), .Q(n820) );
  CLKBU6 U568 ( .A(n822), .Q(n821) );
  CLKBU6 U569 ( .A(n823), .Q(n822) );
  CLKBU6 U570 ( .A(iYa[12]), .Q(n823) );
  CLKBU6 U571 ( .A(n825), .Q(n824) );
  CLKBU6 U572 ( .A(n826), .Q(n825) );
  CLKBU6 U573 ( .A(iXa[13]), .Q(n826) );
  CLKBU6 U574 ( .A(n828), .Q(n827) );
  CLKBU6 U575 ( .A(n829), .Q(n828) );
  CLKBU6 U576 ( .A(n830), .Q(n829) );
  CLKBU6 U577 ( .A(n831), .Q(n830) );
  CLKBU6 U578 ( .A(iYa[13]), .Q(n831) );
  CLKBU6 U579 ( .A(n833), .Q(n832) );
  CLKBU6 U580 ( .A(n834), .Q(n833) );
  CLKBU6 U581 ( .A(iXa[14]), .Q(n834) );
  CLKBU6 U582 ( .A(n836), .Q(n835) );
  CLKBU6 U583 ( .A(n837), .Q(n836) );
  CLKBU6 U584 ( .A(n838), .Q(n837) );
  CLKBU6 U585 ( .A(n839), .Q(n838) );
  CLKBU6 U586 ( .A(iYa[14]), .Q(n839) );
  CLKBU6 U587 ( .A(n841), .Q(n840) );
  CLKBU6 U588 ( .A(n842), .Q(n841) );
  CLKBU6 U589 ( .A(iXa[15]), .Q(n842) );
  CLKBU6 U590 ( .A(n844), .Q(n843) );
  CLKBU6 U591 ( .A(n845), .Q(n844) );
  CLKBU6 U592 ( .A(n846), .Q(n845) );
  CLKBU6 U593 ( .A(n847), .Q(n846) );
  CLKBU6 U594 ( .A(iYa[15]), .Q(n847) );
  CLKBU6 U595 ( .A(n849), .Q(n848) );
  CLKBU6 U596 ( .A(n850), .Q(n849) );
  CLKBU6 U597 ( .A(iXa[16]), .Q(n850) );
  CLKBU6 U598 ( .A(n852), .Q(n851) );
  CLKBU6 U599 ( .A(n853), .Q(n852) );
  CLKBU6 U600 ( .A(n854), .Q(n853) );
  CLKBU6 U601 ( .A(n855), .Q(n854) );
  CLKBU6 U602 ( .A(iYa[16]), .Q(n855) );
  CLKBU6 U603 ( .A(n857), .Q(n856) );
  CLKBU6 U604 ( .A(n858), .Q(n857) );
  CLKBU6 U605 ( .A(iXa[17]), .Q(n858) );
  CLKBU6 U606 ( .A(n860), .Q(n859) );
  CLKBU6 U607 ( .A(n861), .Q(n860) );
  CLKBU6 U608 ( .A(n862), .Q(n861) );
  CLKBU6 U609 ( .A(n863), .Q(n862) );
  CLKBU6 U610 ( .A(iYa[17]), .Q(n863) );
  CLKBU6 U611 ( .A(n865), .Q(n864) );
  CLKBU6 U612 ( .A(n866), .Q(n865) );
  CLKBU6 U613 ( .A(iXa[18]), .Q(n866) );
  CLKBU6 U614 ( .A(n868), .Q(n867) );
  CLKBU6 U615 ( .A(n869), .Q(n868) );
  CLKBU6 U616 ( .A(n870), .Q(n869) );
  CLKBU6 U617 ( .A(n871), .Q(n870) );
  CLKBU6 U618 ( .A(iYa[18]), .Q(n871) );
  CLKBU6 U619 ( .A(n873), .Q(n872) );
  CLKBU6 U620 ( .A(n874), .Q(n873) );
  CLKBU6 U621 ( .A(iXa[19]), .Q(n874) );
  CLKBU6 U622 ( .A(n876), .Q(n875) );
  CLKBU6 U623 ( .A(n877), .Q(n876) );
  CLKBU6 U624 ( .A(n878), .Q(n877) );
  CLKBU6 U625 ( .A(n879), .Q(n878) );
  CLKBU6 U626 ( .A(iYa[19]), .Q(n879) );
  CLKBU6 U627 ( .A(n881), .Q(n880) );
  CLKBU6 U628 ( .A(n882), .Q(n881) );
  CLKBU6 U629 ( .A(iXa[20]), .Q(n882) );
  CLKBU6 U630 ( .A(n884), .Q(n883) );
  CLKBU6 U631 ( .A(n885), .Q(n884) );
  CLKBU6 U632 ( .A(n886), .Q(n885) );
  CLKBU6 U633 ( .A(n887), .Q(n886) );
  CLKBU6 U634 ( .A(iYa[20]), .Q(n887) );
  CLKBU6 U635 ( .A(n889), .Q(n888) );
  CLKBU6 U636 ( .A(n890), .Q(n889) );
  CLKBU6 U637 ( .A(iXa[21]), .Q(n890) );
  CLKBU6 U638 ( .A(n892), .Q(n891) );
  CLKBU6 U639 ( .A(n893), .Q(n892) );
  CLKBU6 U640 ( .A(n894), .Q(n893) );
  CLKBU6 U641 ( .A(n895), .Q(n894) );
  CLKBU6 U642 ( .A(iYa[21]), .Q(n895) );
  CLKBU6 U643 ( .A(n897), .Q(n896) );
  CLKBU6 U644 ( .A(n898), .Q(n897) );
  CLKBU6 U645 ( .A(iXa[22]), .Q(n898) );
  CLKBU6 U646 ( .A(n900), .Q(n899) );
  CLKBU6 U647 ( .A(n901), .Q(n900) );
  CLKBU6 U648 ( .A(n902), .Q(n901) );
  CLKBU6 U649 ( .A(n903), .Q(n902) );
  CLKBU6 U650 ( .A(iYa[22]), .Q(n903) );
  CLKBU6 U651 ( .A(n905), .Q(n904) );
  CLKBU6 U652 ( .A(n906), .Q(n905) );
  CLKBU6 U653 ( .A(iXa[23]), .Q(n906) );
  CLKBU6 U654 ( .A(n908), .Q(n907) );
  CLKBU6 U655 ( .A(n909), .Q(n908) );
  CLKBU6 U656 ( .A(n910), .Q(n909) );
  CLKBU6 U657 ( .A(n911), .Q(n910) );
  CLKBU6 U658 ( .A(iYa[23]), .Q(n911) );
  CLKBU6 U659 ( .A(n913), .Q(n912) );
  CLKBU6 U660 ( .A(n914), .Q(n913) );
  CLKBU6 U661 ( .A(iXa[24]), .Q(n914) );
  CLKBU6 U662 ( .A(n916), .Q(n915) );
  CLKBU6 U663 ( .A(n917), .Q(n916) );
  CLKBU6 U664 ( .A(n918), .Q(n917) );
  CLKBU6 U665 ( .A(n919), .Q(n918) );
  CLKBU6 U666 ( .A(iYa[24]), .Q(n919) );
  CLKBU6 U667 ( .A(n921), .Q(n920) );
  CLKBU6 U668 ( .A(n922), .Q(n921) );
  CLKBU6 U669 ( .A(iXa[25]), .Q(n922) );
  CLKBU6 U670 ( .A(n924), .Q(n923) );
  CLKBU6 U671 ( .A(n925), .Q(n924) );
  CLKBU6 U672 ( .A(n926), .Q(n925) );
  CLKBU6 U673 ( .A(n927), .Q(n926) );
  CLKBU6 U674 ( .A(iYa[25]), .Q(n927) );
  CLKBU6 U675 ( .A(n929), .Q(n928) );
  CLKBU6 U676 ( .A(n930), .Q(n929) );
  CLKBU6 U677 ( .A(iXa[26]), .Q(n930) );
  CLKBU6 U678 ( .A(n932), .Q(n931) );
  CLKBU6 U679 ( .A(n933), .Q(n932) );
  CLKBU6 U680 ( .A(n934), .Q(n933) );
  CLKBU6 U681 ( .A(n935), .Q(n934) );
  CLKBU6 U682 ( .A(iYa[26]), .Q(n935) );
  CLKBU6 U683 ( .A(n937), .Q(n936) );
  CLKBU6 U684 ( .A(n938), .Q(n937) );
  CLKBU6 U685 ( .A(iXa[27]), .Q(n938) );
  CLKBU6 U686 ( .A(n940), .Q(n939) );
  CLKBU6 U687 ( .A(n941), .Q(n940) );
  CLKBU6 U688 ( .A(n942), .Q(n941) );
  CLKBU6 U689 ( .A(n943), .Q(n942) );
  CLKBU6 U690 ( .A(iYa[27]), .Q(n943) );
  CLKBU6 U691 ( .A(n945), .Q(n944) );
  CLKBU6 U692 ( .A(n946), .Q(n945) );
  CLKBU6 U693 ( .A(iXa[28]), .Q(n946) );
  CLKBU6 U694 ( .A(n948), .Q(n947) );
  CLKBU6 U695 ( .A(n949), .Q(n948) );
  CLKBU6 U696 ( .A(n950), .Q(n949) );
  CLKBU6 U697 ( .A(n951), .Q(n950) );
  CLKBU6 U698 ( .A(iYa[28]), .Q(n951) );
  CLKBU6 U699 ( .A(n953), .Q(n952) );
  CLKBU6 U700 ( .A(n954), .Q(n953) );
  CLKBU6 U701 ( .A(iXa[29]), .Q(n954) );
  CLKBU6 U702 ( .A(n956), .Q(n955) );
  CLKBU6 U703 ( .A(n957), .Q(n956) );
  CLKBU6 U704 ( .A(n958), .Q(n957) );
  CLKBU6 U705 ( .A(n959), .Q(n958) );
  CLKBU6 U706 ( .A(iYa[29]), .Q(n959) );
  CLKBU6 U707 ( .A(n961), .Q(n960) );
  CLKBU6 U708 ( .A(n962), .Q(n961) );
  CLKBU6 U709 ( .A(iXa[30]), .Q(n962) );
  CLKBU6 U710 ( .A(n964), .Q(n963) );
  CLKBU6 U711 ( .A(n965), .Q(n964) );
  CLKBU6 U712 ( .A(n966), .Q(n965) );
  CLKBU6 U713 ( .A(n967), .Q(n966) );
  CLKBU6 U714 ( .A(iYa[30]), .Q(n967) );
  CLKBU6 U715 ( .A(n969), .Q(n968) );
  CLKBU6 U716 ( .A(n970), .Q(n969) );
  CLKBU6 U717 ( .A(iXa[31]), .Q(n970) );
  CLKBU6 U718 ( .A(n972), .Q(n971) );
  CLKBU6 U719 ( .A(n973), .Q(n972) );
  CLKBU6 U720 ( .A(n974), .Q(n973) );
  CLKBU6 U721 ( .A(n975), .Q(n974) );
  CLKBU6 U722 ( .A(iYa[31]), .Q(n975) );
  CLKBU6 U723 ( .A(n399), .Q(n976) );
  CLKBU6 U724 ( .A(n976), .Q(n977) );
  CLKBU6 U725 ( .A(n977), .Q(n978) );
  CLKBU6 U726 ( .A(n987), .Q(n986) );
  CLKBU6 U727 ( .A(n987), .Q(n985) );
  CLKBU6 U728 ( .A(n984), .Q(n987) );
  CLKBU6 U729 ( .A(n398), .Q(n984) );
  CLKBU6 U730 ( .A(n269), .Q(n992) );
  CLKBU6 U731 ( .A(n996), .Q(n979) );
  CLKBU6 U732 ( .A(n270), .Q(n988) );
  CLKBU6 U733 ( .A(n270), .Q(n989) );
  CLKBU6 U734 ( .A(n270), .Q(n990) );
  CLKBU6 U735 ( .A(n270), .Q(n991) );
  CLKBU6 U736 ( .A(n269), .Q(n993) );
  CLKBU6 U737 ( .A(n269), .Q(n994) );
  CLKBU6 U738 ( .A(n996), .Q(n980) );
  NAND22 U739 ( .A(n995), .B(n265), .Q(n269) );
  CLKBU6 U740 ( .A(n998), .Q(n982) );
  NOR22 U741 ( .A(n397), .B(n992), .Q(n270) );
  CLKBU6 U742 ( .A(n998), .Q(n983) );
  AOI2111 U743 ( .A(n262), .B(iEn), .C(n982), .D(n979), .Q(n399) );
  NAND22 U744 ( .A(R_STATE__0_), .B(n262), .Q(n266) );
  NAND22 U745 ( .A(R_STATE__1_), .B(n264), .Q(n265) );
  NAND22 U746 ( .A(n329), .B(n330), .Q(n430) );
  AOI221 U747 ( .A(n728), .B(n990), .C(R_YA__1_), .D(n998), .Q(n329) );
  NAND22 U748 ( .A(n321), .B(n322), .Q(n426) );
  NAND22 U749 ( .A(R_XA__5_), .B(n993), .Q(n322) );
  AOI221 U750 ( .A(n760), .B(n990), .C(R_YA__5_), .D(n983), .Q(n321) );
  NAND22 U751 ( .A(n317), .B(n318), .Q(n424) );
  NAND22 U752 ( .A(R_XA__7_), .B(n994), .Q(n318) );
  AOI221 U753 ( .A(n776), .B(n991), .C(R_YA__7_), .D(n998), .Q(n317) );
  NAND22 U754 ( .A(n313), .B(n314), .Q(n422) );
  NAND22 U755 ( .A(R_XA__9_), .B(n994), .Q(n314) );
  AOI221 U756 ( .A(n792), .B(n988), .C(R_YA__9_), .D(n983), .Q(n313) );
  NAND22 U757 ( .A(n309), .B(n310), .Q(n420) );
  NAND22 U758 ( .A(R_XA__11_), .B(n994), .Q(n310) );
  AOI221 U759 ( .A(n808), .B(n989), .C(R_YA__11_), .D(n998), .Q(n309) );
  NAND22 U760 ( .A(n305), .B(n306), .Q(n418) );
  NAND22 U761 ( .A(R_XA__13_), .B(n994), .Q(n306) );
  AOI221 U762 ( .A(n824), .B(n990), .C(R_YA__13_), .D(n983), .Q(n305) );
  NAND22 U763 ( .A(n301), .B(n302), .Q(n416) );
  NAND22 U764 ( .A(R_XA__15_), .B(n994), .Q(n302) );
  AOI221 U765 ( .A(n840), .B(n991), .C(R_YA__15_), .D(n982), .Q(n301) );
  NAND22 U766 ( .A(n297), .B(n298), .Q(n414) );
  NAND22 U767 ( .A(R_XA__17_), .B(n994), .Q(n298) );
  AOI221 U768 ( .A(n856), .B(n988), .C(R_YA__17_), .D(n982), .Q(n297) );
  NAND22 U769 ( .A(n293), .B(n294), .Q(n412) );
  NAND22 U770 ( .A(R_XA__19_), .B(n994), .Q(n294) );
  AOI221 U771 ( .A(n872), .B(n989), .C(R_YA__19_), .D(n982), .Q(n293) );
  NAND22 U772 ( .A(n289), .B(n290), .Q(n410) );
  NAND22 U773 ( .A(R_XA__21_), .B(n994), .Q(n290) );
  AOI221 U774 ( .A(n888), .B(n991), .C(R_YA__21_), .D(n982), .Q(n289) );
  NAND22 U775 ( .A(n285), .B(n286), .Q(n408) );
  NAND22 U776 ( .A(R_XA__23_), .B(n994), .Q(n286) );
  AOI221 U777 ( .A(n904), .B(n991), .C(R_YA__23_), .D(n982), .Q(n285) );
  NAND22 U778 ( .A(n281), .B(n282), .Q(n406) );
  NAND22 U779 ( .A(R_XA__25_), .B(n993), .Q(n282) );
  AOI221 U780 ( .A(n920), .B(n991), .C(R_YA__25_), .D(n982), .Q(n281) );
  NAND22 U781 ( .A(n277), .B(n278), .Q(n404) );
  NAND22 U782 ( .A(R_XA__27_), .B(n993), .Q(n278) );
  AOI221 U783 ( .A(n936), .B(n991), .C(R_YA__27_), .D(n982), .Q(n277) );
  NAND22 U784 ( .A(n273), .B(n274), .Q(n402) );
  NAND22 U785 ( .A(R_XA__29_), .B(n994), .Q(n274) );
  AOI221 U786 ( .A(n952), .B(n991), .C(R_YA__29_), .D(n982), .Q(n273) );
  NAND22 U787 ( .A(n267), .B(n268), .Q(n400) );
  NAND22 U788 ( .A(R_XA__31_), .B(n993), .Q(n268) );
  AOI221 U789 ( .A(n968), .B(n991), .C(R_YA__31_), .D(n983), .Q(n267) );
  NAND22 U790 ( .A(n325), .B(n326), .Q(n428) );
  NAND22 U791 ( .A(R_XA__3_), .B(n993), .Q(n326) );
  AOI221 U792 ( .A(n744), .B(n990), .C(R_YA__3_), .D(n998), .Q(n325) );
  NAND22 U793 ( .A(n327), .B(n328), .Q(n429) );
  NAND22 U794 ( .A(R_XA__2_), .B(n994), .Q(n328) );
  AOI221 U795 ( .A(n736), .B(n990), .C(R_YA__2_), .D(n983), .Q(n327) );
  NAND22 U796 ( .A(n331), .B(n332), .Q(n431) );
  NAND22 U797 ( .A(R_XA__0_), .B(n993), .Q(n332) );
  AOI221 U798 ( .A(n720), .B(n990), .C(R_YA__0_), .D(n998), .Q(n331) );
  NAND22 U799 ( .A(n395), .B(n396), .Q(n463) );
  NAND22 U800 ( .A(R_XB__0_), .B(n992), .Q(n396) );
  AOI221 U801 ( .A(n464), .B(n988), .C(R_YB__0_), .D(n983), .Q(n395) );
  NAND22 U802 ( .A(n393), .B(n394), .Q(n462) );
  NAND22 U803 ( .A(R_XB__1_), .B(n992), .Q(n394) );
  AOI221 U804 ( .A(n472), .B(n988), .C(R_YB__1_), .D(n983), .Q(n393) );
  NAND22 U805 ( .A(n391), .B(n392), .Q(n461) );
  NAND22 U806 ( .A(R_XB__2_), .B(n992), .Q(n392) );
  AOI221 U807 ( .A(n480), .B(n988), .C(R_YB__2_), .D(n983), .Q(n391) );
  NAND22 U808 ( .A(n389), .B(n390), .Q(n460) );
  NAND22 U809 ( .A(R_XB__3_), .B(n992), .Q(n390) );
  AOI221 U810 ( .A(n488), .B(n988), .C(R_YB__3_), .D(n983), .Q(n389) );
  NAND22 U811 ( .A(n387), .B(n388), .Q(n459) );
  NAND22 U812 ( .A(R_XB__4_), .B(n992), .Q(n388) );
  AOI221 U813 ( .A(n496), .B(n988), .C(R_YB__4_), .D(n983), .Q(n387) );
  NAND22 U814 ( .A(n385), .B(n386), .Q(n458) );
  NAND22 U815 ( .A(R_XB__5_), .B(n992), .Q(n386) );
  AOI221 U816 ( .A(n504), .B(n988), .C(R_YB__5_), .D(n983), .Q(n385) );
  NAND22 U817 ( .A(n383), .B(n384), .Q(n457) );
  NAND22 U818 ( .A(R_XB__6_), .B(n992), .Q(n384) );
  AOI221 U819 ( .A(n512), .B(n988), .C(R_YB__6_), .D(n983), .Q(n383) );
  NAND22 U820 ( .A(n381), .B(n382), .Q(n456) );
  NAND22 U821 ( .A(R_XB__7_), .B(n992), .Q(n382) );
  AOI221 U822 ( .A(n520), .B(n988), .C(R_YB__7_), .D(n983), .Q(n381) );
  NAND22 U823 ( .A(n379), .B(n380), .Q(n455) );
  NAND22 U824 ( .A(R_XB__8_), .B(n992), .Q(n380) );
  AOI221 U825 ( .A(n528), .B(n988), .C(R_YB__8_), .D(n983), .Q(n379) );
  NAND22 U826 ( .A(n377), .B(n378), .Q(n454) );
  NAND22 U827 ( .A(R_XB__9_), .B(n992), .Q(n378) );
  AOI221 U828 ( .A(n536), .B(n988), .C(R_YB__9_), .D(n983), .Q(n377) );
  NAND22 U829 ( .A(n375), .B(n376), .Q(n453) );
  NAND22 U830 ( .A(R_XB__10_), .B(n992), .Q(n376) );
  AOI221 U831 ( .A(n544), .B(n988), .C(R_YB__10_), .D(n983), .Q(n375) );
  NAND22 U832 ( .A(n373), .B(n374), .Q(n452) );
  NAND22 U833 ( .A(R_XB__11_), .B(n992), .Q(n374) );
  AOI221 U834 ( .A(n552), .B(n988), .C(R_YB__11_), .D(n983), .Q(n373) );
  NAND22 U835 ( .A(n371), .B(n372), .Q(n451) );
  NAND22 U836 ( .A(R_XB__12_), .B(n993), .Q(n372) );
  AOI221 U837 ( .A(n560), .B(n988), .C(R_YB__12_), .D(n983), .Q(n371) );
  NAND22 U838 ( .A(n369), .B(n370), .Q(n450) );
  NAND22 U839 ( .A(R_XB__13_), .B(n993), .Q(n370) );
  AOI221 U840 ( .A(n568), .B(n989), .C(R_YB__13_), .D(n983), .Q(n369) );
  NAND22 U841 ( .A(n367), .B(n368), .Q(n449) );
  NAND22 U842 ( .A(R_XB__14_), .B(n993), .Q(n368) );
  AOI221 U843 ( .A(n576), .B(n989), .C(R_YB__14_), .D(n983), .Q(n367) );
  NAND22 U844 ( .A(n365), .B(n366), .Q(n448) );
  NAND22 U845 ( .A(R_XB__15_), .B(n993), .Q(n366) );
  AOI221 U846 ( .A(n584), .B(n989), .C(R_YB__15_), .D(n983), .Q(n365) );
  NAND22 U847 ( .A(n363), .B(n364), .Q(n447) );
  NAND22 U848 ( .A(R_XB__16_), .B(n993), .Q(n364) );
  AOI221 U849 ( .A(n592), .B(n989), .C(R_YB__16_), .D(n983), .Q(n363) );
  NAND22 U850 ( .A(n361), .B(n362), .Q(n446) );
  NAND22 U851 ( .A(R_XB__17_), .B(n993), .Q(n362) );
  AOI221 U852 ( .A(n600), .B(n989), .C(R_YB__17_), .D(n983), .Q(n361) );
  NAND22 U853 ( .A(n359), .B(n360), .Q(n445) );
  NAND22 U854 ( .A(R_XB__18_), .B(n993), .Q(n360) );
  AOI221 U855 ( .A(n608), .B(n989), .C(R_YB__18_), .D(n983), .Q(n359) );
  NAND22 U856 ( .A(n357), .B(n358), .Q(n444) );
  NAND22 U857 ( .A(R_XB__19_), .B(n993), .Q(n358) );
  AOI221 U858 ( .A(n616), .B(n989), .C(R_YB__19_), .D(n983), .Q(n357) );
  NAND22 U859 ( .A(n355), .B(n356), .Q(n443) );
  NAND22 U860 ( .A(R_XB__20_), .B(n993), .Q(n356) );
  AOI221 U861 ( .A(n624), .B(n989), .C(R_YB__20_), .D(n983), .Q(n355) );
  NAND22 U862 ( .A(n353), .B(n354), .Q(n442) );
  NAND22 U863 ( .A(R_XB__21_), .B(n993), .Q(n354) );
  AOI221 U864 ( .A(n632), .B(n989), .C(R_YB__21_), .D(n983), .Q(n353) );
  NAND22 U865 ( .A(n351), .B(n352), .Q(n441) );
  NAND22 U866 ( .A(R_XB__22_), .B(n993), .Q(n352) );
  AOI221 U867 ( .A(n640), .B(n989), .C(R_YB__22_), .D(n983), .Q(n351) );
  NAND22 U868 ( .A(n349), .B(n350), .Q(n440) );
  NAND22 U869 ( .A(R_XB__23_), .B(n993), .Q(n350) );
  AOI221 U870 ( .A(n648), .B(n989), .C(R_YB__23_), .D(n983), .Q(n349) );
  NAND22 U871 ( .A(n347), .B(n348), .Q(n439) );
  NAND22 U872 ( .A(R_XB__24_), .B(n993), .Q(n348) );
  AOI221 U873 ( .A(n656), .B(n989), .C(R_YB__24_), .D(n983), .Q(n347) );
  NAND22 U874 ( .A(n345), .B(n346), .Q(n438) );
  NAND22 U875 ( .A(R_XB__25_), .B(n993), .Q(n346) );
  AOI221 U876 ( .A(n664), .B(n989), .C(R_YB__25_), .D(n983), .Q(n345) );
  NAND22 U877 ( .A(n315), .B(n316), .Q(n423) );
  NAND22 U878 ( .A(R_XA__8_), .B(n994), .Q(n316) );
  AOI221 U879 ( .A(n784), .B(n990), .C(R_YA__8_), .D(n983), .Q(n315) );
  NAND22 U880 ( .A(n311), .B(n312), .Q(n421) );
  NAND22 U881 ( .A(R_XA__10_), .B(n994), .Q(n312) );
  AOI221 U882 ( .A(n800), .B(n991), .C(R_YA__10_), .D(n998), .Q(n311) );
  NAND22 U883 ( .A(n307), .B(n308), .Q(n419) );
  NAND22 U884 ( .A(R_XA__12_), .B(n994), .Q(n308) );
  AOI221 U885 ( .A(n816), .B(n270), .C(R_YA__12_), .D(n998), .Q(n307) );
  NAND22 U886 ( .A(n303), .B(n304), .Q(n417) );
  NAND22 U887 ( .A(R_XA__14_), .B(n994), .Q(n304) );
  AOI221 U888 ( .A(n832), .B(n270), .C(R_YA__14_), .D(n983), .Q(n303) );
  NAND22 U889 ( .A(n299), .B(n300), .Q(n415) );
  NAND22 U890 ( .A(R_XA__16_), .B(n994), .Q(n300) );
  AOI221 U891 ( .A(n848), .B(n270), .C(R_YA__16_), .D(n982), .Q(n299) );
  NAND22 U892 ( .A(n295), .B(n296), .Q(n413) );
  NAND22 U893 ( .A(R_XA__18_), .B(n994), .Q(n296) );
  AOI221 U894 ( .A(n864), .B(n270), .C(R_YA__18_), .D(n982), .Q(n295) );
  NAND22 U895 ( .A(n291), .B(n292), .Q(n411) );
  NAND22 U896 ( .A(R_XA__20_), .B(n994), .Q(n292) );
  AOI221 U897 ( .A(n880), .B(n991), .C(R_YA__20_), .D(n982), .Q(n291) );
  NAND22 U898 ( .A(n343), .B(n344), .Q(n437) );
  NAND22 U899 ( .A(R_XB__26_), .B(n994), .Q(n344) );
  AOI221 U900 ( .A(n672), .B(n990), .C(R_YB__26_), .D(n983), .Q(n343) );
  NAND22 U901 ( .A(n341), .B(n342), .Q(n436) );
  NAND22 U902 ( .A(R_XB__27_), .B(n993), .Q(n342) );
  AOI221 U903 ( .A(n680), .B(n990), .C(R_YB__27_), .D(n983), .Q(n341) );
  NAND22 U904 ( .A(n339), .B(n340), .Q(n435) );
  NAND22 U905 ( .A(R_XB__28_), .B(n994), .Q(n340) );
  AOI221 U906 ( .A(n688), .B(n990), .C(R_YB__28_), .D(n983), .Q(n339) );
  NAND22 U907 ( .A(n337), .B(n338), .Q(n434) );
  NAND22 U908 ( .A(R_XB__29_), .B(n993), .Q(n338) );
  AOI221 U909 ( .A(n696), .B(n990), .C(R_YB__29_), .D(n983), .Q(n337) );
  NAND22 U910 ( .A(n335), .B(n336), .Q(n433) );
  NAND22 U911 ( .A(R_XB__30_), .B(n994), .Q(n336) );
  AOI221 U912 ( .A(n704), .B(n990), .C(R_YB__30_), .D(n983), .Q(n335) );
  NAND22 U913 ( .A(n333), .B(n334), .Q(n432) );
  NAND22 U914 ( .A(R_XB__31_), .B(n993), .Q(n334) );
  AOI221 U915 ( .A(n712), .B(n990), .C(R_YB__31_), .D(n998), .Q(n333) );
  NAND22 U916 ( .A(n323), .B(n324), .Q(n427) );
  NAND22 U917 ( .A(R_XA__4_), .B(n994), .Q(n324) );
  AOI221 U918 ( .A(n752), .B(n990), .C(R_YA__4_), .D(n983), .Q(n323) );
  NAND22 U919 ( .A(n319), .B(n320), .Q(n425) );
  NAND22 U920 ( .A(R_XA__6_), .B(n993), .Q(n320) );
  AOI221 U921 ( .A(n768), .B(n990), .C(R_YA__6_), .D(n982), .Q(n319) );
  NAND22 U922 ( .A(n287), .B(n288), .Q(n409) );
  NAND22 U923 ( .A(R_XA__22_), .B(n993), .Q(n288) );
  AOI221 U924 ( .A(n896), .B(n991), .C(R_YA__22_), .D(n982), .Q(n287) );
  NAND22 U925 ( .A(n283), .B(n284), .Q(n407) );
  NAND22 U926 ( .A(R_XA__24_), .B(n994), .Q(n284) );
  AOI221 U927 ( .A(n912), .B(n991), .C(R_YA__24_), .D(n998), .Q(n283) );
  NAND22 U928 ( .A(n279), .B(n280), .Q(n405) );
  NAND22 U929 ( .A(R_XA__26_), .B(n993), .Q(n280) );
  AOI221 U930 ( .A(n928), .B(n991), .C(R_YA__26_), .D(n982), .Q(n279) );
  NAND22 U931 ( .A(n275), .B(n276), .Q(n403) );
  NAND22 U932 ( .A(R_XA__28_), .B(n994), .Q(n276) );
  AOI221 U933 ( .A(n944), .B(n991), .C(R_YA__28_), .D(n982), .Q(n275) );
  NAND22 U934 ( .A(n271), .B(n272), .Q(n401) );
  NAND22 U935 ( .A(R_XA__30_), .B(n994), .Q(n272) );
  AOI221 U936 ( .A(n960), .B(n991), .C(R_YA__30_), .D(n982), .Q(n271) );
  NAND22 U937 ( .A(n264), .B(n262), .Q(n397) );
  NAND22 U938 ( .A(R_XA__1_), .B(n994), .Q(n330) );
  CLKIN6 U939 ( .A(n978), .Q(n995) );
  CLKIN6 U940 ( .A(n266), .Q(n998) );
endmodule

